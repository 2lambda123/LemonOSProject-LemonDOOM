ELF          >    @     @       0l!         @ 8  @ # "       @       @ @     @ @                              X      X@     X@                                          @       @     ,Y     ,Y                   0Y     0Yd     0Yd     �:     `                   XY     XYd     XYd     �      �             /lib/ld64.so.1  %   -   +   #   *                                !           )             (   $         '   ,                          %                                                                                                                                                    
                  &   "       	                              �     ��e            .                      �                      �                      6                      �                      '                      M                      �                                                                   u                      �                      �                      `                      �                                           n                                           T                      �                                           �                      /   	 @            �                      	                      �                                           �                      }                                           ?                                           5                                            �                      #                     �                      �                                           �                      (                     �                      �                       libc.so putchar strcpy tolower system malloc remove vsnprintf __mlibc_errno fflush strncasecmp __mlibc_entry rename strrchr calloc atof fseek strstr strncmp strncpy strcasecmp realloc sscanf fread strdup fopen ftell fclose strcmp stderr fwrite exit atoi toupper strchr fputs mkdir vfprintf free memcpy _start   �Zd                    ��e                   �Zd                    [d                   [d                   [d                   [d                    [d                   ([d                   0[d        	           8[d        
           @[d                   H[d                   P[d                   X[d                   `[d                   h[d                   p[d                   x[d                   �[d                   �[d                   �[d                   �[d                   �[d                   �[d                   �[d                   �[d                   �[d                   �[d                   �[d                   �[d                   �[d        !           �[d        "           �[d        #           �[d        $            \d        %           \d        &           \d        '           \d        (            \d        )           (\d        *           0\d        +           8\d        ,           ��  �&> �     �5�N$ �%�N$ @ �%�N$ h    ������%�N$ h   ������%�N$ h   ������%�N$ h   �����%�N$ h   �����%zN$ h   �����%rN$ h   �����%jN$ h   �p����%bN$ h   �`����%ZN$ h	   �P����%RN$ h
   �@����%JN$ h   �0����%BN$ h   � ����%:N$ h   �����%2N$ h   � ����%*N$ h   ������%"N$ h   ������%N$ h   ������%N$ h   ������%
N$ h   �����%N$ h   �����%�M$ h   �����%�M$ h   �����%�M$ h   �p����%�M$ h   �`����%�M$ h   �P����%�M$ h   �@����%�M$ h   �0����%�M$ h   � ����%�M$ h   �����%�M$ h   � ����%�M$ h   ������%�M$ h    ������%�M$ h!   ������%�M$ h"   ������%�M$ h#   �����%�M$ h$   �����%zM$ h%   �����%rM$ h&   �����%jM$ h'   �p����%bM$ h(   �`���PH�5@5& �=25& �A  ��JB ����1��� �W+  1�Z�H�h&     �H���@ �����f.�     ��ؓe H=ؓe t�    H��t	�ؓe ��f��ff.�     @ �ؓe H��ؓe H��H��H��?H�H��t�    H��t�ؓe ���ff.�     @ �=Y�%  uwUH�W�% H��ATA�HYd S�PYd H��HYd H��H��H9�s%f.�     H��H��% A��H��% H9�r��0����    H��t
��C ����[A\��% ]��ff.�     @ �    H��tU� �e ��C H�����]����D  �����ATI��US�_�o++ou����������F��t�"����;�  A�D$��u�  ���x�����	�މ���  []A�$A\Ë��% �=0�% S�   �5��% ������% �΄% ���Մ% �ƈ  �=��% �5x�% ���% ��謈  �5��% �����% ���% ���)Ɖș�5��% �����% [)w�% щ{�% ��k�% �i�% Ëj�% �(�% �Z�% ��% �B�% ��% �2�% ��% �R�5�% ���% �=KK$  �5�% ��% u�ۃ% ��% �˃% ��% �1H���% �   L� ����A�P)ȉ�% ���A�P)΃% �̃% �=��% ��% ������% ���% 讇  �   �Ɖ�J$ 蜇  �B�% XËz�% �   Hc=n�% ���u�% ����e �T�% ����
   V�% ��Ĕe �G����7�% �� �% ���1�E1ɺ  �ATD�%�L& E1�E1�UH�-;M& ��������% ���A�����ւ%   ��Ђ%   �S1�A9�~6�L� D9�|9�~��A��A�ȳ�L�9�|9�~��A����A�H���ń�tD���% E��t�=|�% E��t�5u�% E��t�b�% �=��% �5Z�% �P�% +5V�% +L�% ���7�% �^�  �=��% �5&�% �����H�  �=j�% �    9�O������% �*�  []��% A\Ë5%�% �#�% ��	�t�I$     ���% ����=߁% A�   5�% �5݁% Ӂ% ���ˁ% �A�����% �9�
���% 9�})��% �5��% A�   ��A���q�% �9�
�m�% 9�})y�% �w�% 5m�% �5_�% ��[�% �R�=��% H��& �5��% ��%    ��% �����H�P�% �>�%     �D�%     H�!�%     ��%    ��%    ��  �=�% �5��% �ր% ���Є  A�����% Hc�!& �<��9f  uH�a�% �;f 1҃<��9f  Hc�tHi�H  H�;f H�>�% �	H��H��u�H�,�% D�m�% �   H�0D�Й���V)�D�ȉa�% ����V)O�% �3����H�% �p\d D��% ��% �,�% D��% ��% X�{� S1�H���ٺ�JB �	   1�H�|$�����   H�|$� H�� �e H��H��
u�H��[�S1�H���ٺ�JB �	   1�H�|$���o���H�|$� ��
u�H��[�1�����e ����H��H��
u��r~%     �R��%     ��%     ��% @  ��% �   ���������=% �3�  �B�  ;% �VF$ ~��~% �HF$ �5BF$ �   ��  ��~% X�P�.����P\d ��}%     �P� ��E$    Z�R�=�E$  u�������E$     �*& 9=E$ u�"& 9+E$ t�+�����)& �E$ ��!& �E$ �-���X�l���P�5V~% �   �5�E$ �v�  �~% Z�Z���P�5/~% �   �5xE$ �S�  ��}% Z�7���UH��SQ�=�|%  �u21ۅ��6  ��9% 9G�'  �.����   ��#&     �  ����  �G9�9% u!1ۃ=E$  �6  �5�}% �   ���  �)9^9% u,1ۃ=�D$  �  �5_}% �   藁  �؉�}% ��  969% u!1ۃ=�D$  ��  �5+}% �   �c�  �)9	9% u,1ۃ=~D$  ��  �5}% �   �:�  �؉T}% �  9�8% u�1}% ��  �#}%  �m  9�8% u�}%  �}% ��  �L  98% u��{%     ��"&    ������&  9U8% u.��{% 1҅���{% u�A����#�����   �c�����   98% uF��C$ 1��;|% ���������C$ H�|% uHǀ�   �JB �   Hǀ�   �JB �   9�7% u6�}|% 1������p|% H��{% uHǀ�   �JB �qHǀ�   KB �d9�7% u;D��z% �KB �KB 1��   ���e �5�  H��{% Hǀ�   ��e �@����!1�9>7% u����H�`{% Hǀ�    KB �   �=�&  ��   �u��\d �]t  ����   ��{% �   �������{% �y1���uu�G9�6% u�vB$ ��u^�X{%     �T9�6% t�9�6% u�PB$ ��u8�6{%     �.9�6% t�9�6% t9�6% u�{%    ��z%    1ۉ�Z[]�V�5�z% �=B$ ��~  �   �Ɖ�A$ ��~  �rz% ��A$ ;�z% }Y�%���;xz% ~Z�:���X����H�;z% H� �x9=?z% u�@98z% ��   USP�5�A$ �z% �T~  �޻   f1����C~  �5oA$ �-�y% ���-z% ���)�H��y% �+z% H� �x�~  ��f1����~  ����y% �����y% �y% ��y% )����y% ��y% ��y% H��y% H� H�@H��y% Z[]�Ë�y% ;�x% ~?Hc~x% �J��`KB �nx% ��y% ��u
�Yx%     �   ��H��)щJx% Ã=
x%  t<Q��y% �=�@$  t������=Uy%    t�^����Ty% Ry% tZ����X�Ë]y% �Ry% ��H�==y% Hc���AUATUS�   Q�G��x% 9�1�;�x% �����W�   9�|1�;�x% ������t1��  ���x% 9�}���;�x% ~��D�GD9�~���D;�x% ~��!�u�H��)ʋ5�?$ I�����n|  �5�?$ A�|$���x% +=^x% �E D�-�x% �E|  �5q?$ A�|$��+=?x% A)�D-ix% D�m�|  �5J?$ A�|$��Px% +=x% �ED�-4x% ��{  �U�   ��A)ŋ#x% D�E��x1�;	x% @�����U ��y���;�w% |����x;�w% �   M���   �E��y���;�w% |���������D��w% D��w% E�Q�E�X���	��  ����E�@��t!�M �ED�e)�A��D+e�A���1��   @��t$D�e�M �ED��D+e)�D)��A���D���W����t'�M D�eD�ҋE)�D)��U)ʉљ��D��D��)����t D�e�U D�mD��+E��A)ՙA��D����9�u.�M �   �E��x1�A9�@������y���5A9�0���+�M�   �E��x1�A9�������y���A9�����������|����   Z[]A\A]�D�E��x7D�bv% E9�}+�O��x$D�Kv% D9�}�WA9�~��x�GA9�~��y"��t% H�=t% �2KB �B��t% 1������D)�)�AUA�   A��A��ATL�%�u% A��A��UD1�D1�SD)�D)�A��A����, 9�~2�ؙA����)�D����D�Hc�A�4D9GtJ��xD�)�E���ډ�A����E��E��)�D����F� Mc�C�49Ot��xE�)�D��D���[]A\A]�S�󾀔e ������t�޿��e [�����[�ATU��SH����t% ��+q?& �˩�� t�  � ���)�ˋ�t% �t% A�̉D$�t% �D$D9�}��H��$�\$��  � �z������t% ��+?& �˩�� t�  � ���)�ˋxt% ^t% A�̉$Vt% �D$D9�}��H��\$�\$��  � ������H��[]A\�S1�9�>& ��   Hk�XH�>& �5Zt% H��
�R��r% H�P��r% �
�R��r% ��r% �P��u��tm���   H�H@H��tf�x'u��   �d�� t��s% ���   �QH�@8�899t��s% �p@�<�@9At��s% ���   �&��t,��s% �p`�H�s% �xH t��u�c   �p�e �.���H������[���H��i% AVAUI��ATUH��S�Ӌ?�4��w  D�4���B A�} A��D���w  �} D��A)���v  A�} A��H��i% �4���v  [A�E�u D�e ]A\A]A^�AWE��AVE��AUE1�ATA��U��SH��H��(�t$D;l$��   �3�C�t$�D$��t���v  �t$��D$�wv  �D$E��tH�t$D��H�|$�����D$`�sD$�CDt$�t$�D$��t���6v  �t$��D$�'v  �D$E��tH�t$H�|$D�������D��H�|$�D$`A��Dt$H��D$������=���H��([]A\A]A^A_�USS�=�&  uSH�zq% �=r%  H� �PD�H�H8tA��   AS�   ��]d R1��A��   AR�   ��^d R1�����_AX�r��;f 1ۃ=�&  t�=�&  u	H9-q% u?���9f  t6�}@ A��   uD��@KB H�E �   ��^d �H8D�HR1ҋ@P�M���Y^H��H��H  H��u�X[]�ATA��U1�S9-�;& ~NH��H��H�;& H�X`H��t2�K8D�KP�   �C�   � ]d D��p% PE������ZH�[(Y��H���[]A\�ATE1�USA��$��e ���t�5�7$ +=�p% �yt  �5�7$ A��$Ĕe ��+=lp% �p% �Ë-�p% �Ot  9�p% <����p% )ŋtp% �t ��9�| 9��[p% ��9�|I��$ �e ���q� I��I��P�f���[]A\Ë,p% �   ���"p% ���H�p% H�@�<Ã=rn%  tjR1������=p%  t
�h   �����~���������=�o% u�   �p   �����`   �����������o% ��o% �5�o% �=�o% X�� �Hc�o% H��Hk����@�e �O��P�e �@   �����o% Ë�o% 1�;�o% tHc����@   �Hk���H��@�e �eo% H���I���1�I��L���H��H��J�	L���1�H��J�<	H9�wH)�A�|�/uPI�<�����Z�������Ë0t% ��Hc���H��`�e �XB �t% �AUATI��UL��SV艌  ����   ����1�9�s% Hc�~lL�,�`�e L��L���S�����t L���P�  ��tH�<�`�e Y[]A\A]����H�<�`�e 1�L��1��(�B H����  H��H����  ��uH�������1�ZH��[]A\A]�SH���R���H��HD�[�AWAVI���   AUATUSH���|$��NB ��e  ����   H�& H�H�\�H������I��H��uH�޿�NB 1��a  �/   L��M������H��tL�`1ۋ��PB �D$��sH���PB L���Z�����tH��H��P  uѽ	   A�.��   ��NB E1�������d���D9%�r% ��   J�,�`�e 1�D���PB �D$D����   L���PB H��L���������tH���؊  ��tH������I���W��XB H��������u
L��������1�L��(�B H��1��}�  I��H�ƿ�NB 1��N���L���~�  ��u
L���
����
M��tE�>�H��H��P  �J���E1�I��M���$����E1�H��L��[]A\A]A^A_�AUA���x   ATU1�S1�Q�����I�ċ��PB A��s!H���PB �a���H��tHc�H���PB ��I��H��H��P  u�Hc�L��I��    Z[]A\A]�1�Hk�9��PB uH���PB �H��H��u�
OB ú�PB 1�9zu9ruH�Hk�H���PB ���H����uݸ
OB ú�PB 1�9zu��uH�Hk�H���PB �9rt���H����uظOB �Ë�i% ��t%1�1��   ��u1Ƀ<���e  ��H��H��u߃=�i%  �   D��Q��b  �=}5$  ��t�o& �   ����k�#��  ���Z�USH���H& �-N& �@ H��t% 1��H��t% 1��R1Ƀ=i%  ��   �؋5�t% �5$ �����)ǅ�t��h% ��u���
1Ƀ����TH�Lt% W�H��$�P�It% ��   $����7t% ���   �*t% Hc�HiҠ   ǂ`�e    )���e H����[]Ã=�s%  uVUSR�������=z& ��+n& �h& ��s% 9�|��s%     ��1�)��)ȉ�s% ��������t��9�u�X[]��H��SD�h% H	�uE��t��QB 1���\  ��QB [�:���1�A��   D��D�ds% 	�t=D��H��LcəH��A����Hc�Hk�
Hk�(L�H��)���e I�D ����e H��H��u�A��[D�s% �P�
�����=� & �� & ZË�r% H�G<   �G,    �GDH�      H��V3$     �P &    �S�   H����*@ �E[  �C@[�Zr% 1��AWAVAUATUSR�G`  D�- r% ��= & �=r%  �ŉ
r% t������b������% D�%[r% �D���=��% )Ã=�2$  ��   ��C�D)�9�~���9�O˅ɻ   Oك=�f%  �	  ��q% 1�����q% �<���e  t	��u��   H��H��u���   ��q% A9��\�% ��;cq% D�%\q% ���҉�p�e �=Pq%  ��   �=Gq%  ��   �=>q%  ��   �=5q%  tz�uq%    �n�۸   N��b���% ��=��% �D9���   �L������% D�%Eq% ��=��% D9�~�RB 1��Z  ��^  ��=��% )���2  �   �_  �������u�뫋|�% ���D9�~�/RB 1��WZ  A(A(NL��H��H��p% )�p% )�p% �P�;�% L��1Ҁ��e  ƀ�e  yƀ�e  ��H����u�A�ǋ�% D9���{����˃����   �0�������   ���% ��   ��=��% ���Hc�Li�   �=�d%  I����e uFǅ�       ǅ�       ǅ�       ǅ�       ǅ�       ǅ�       ǅ�       M��`�e E1��T���X[]A\A]A^A_�H�=�o% ËKd% 1��& �& u�	& �& 	�% ����Ã=/0$  tA�=��%  t8�=��%  u/R�>RB ��]  ���   �LRB �� H���U  1��Z���X�Ã=��%  t�S����H��H��tH���Nx  ��u�H����.  ��[�U��jd S1�H����h  �.� �T  �W  �a  �e  �`f  �g  �   �h  ��Ze �SRB H�g   i   H�=& H�b   r   H�4& �_  �t�e �eRB �_  �p�e �pRB �_  ��Ze �}RB �_  ��Ze ��RB �v_  ���e ��RB �g_  �l�e ��RB �X_  ��ed ��RB �I_  ��ed ��RB �:_  �d`d ��RB �+_  �ٺ�RB �   1�H�|$���\�  H��H�|$H��� _  ��
u�H��[]��W�% y
�G�%    �PH�=~�% �   �s� 1�1�YH���� ATUSH����	& ���3  �=��&  t��k �%.$ �������%    �.$ 9�& t��   �@  1�1��$  �   �=�&  u�=��%  t4�=N  ��& ����   ��t����   ����   �B����   �=��%  ty�=�a%  t�#������& �ޅ�u=�   t1��=�%  @�ƃ=�%  t�=�&  �   D�1�=�   @���϶ 1��=@�& �   ���ϼ% ��P� ��  �$� �=�&  uE�=a%  t�=�%  t\�:M  �,�=��%  tLHc=& Hi�H  H���;f �n �=�&  tċ�& 9�,$ t��t��RB �   ��� H���� �=~&  uq�=�,$  u�=�`%  t�]��%     �b �=R&  t��C�=T�& @  t7�& �% u	�=�%  u��%    �	�=ܻ%  t�fd �ϻ% �=T�%  t�=�& �s� ��& �=~&  ���% �j& ���% �& ���% ��& ��+$ ��+$ tL�=�_%  �   u	���& �h�   ��RB ��� �   H�Ƌ��& ��D���H�����& ���T� �.q  �������uH��[]A\�z� ��   �@  1�1��!  �X  �X��X  �   A����A)�D�L$�X  D�L$E��~�A��   �@  1�1��   ���!  A���� �p  �� E��t�H��[]A\�P�=�%  t!�=�& t�l& >& t�SB �
����=+&  t�S:  �B�%    ����H�=��% �7� �7� ��/@ �.� ��� �%� �M� �Ah ������=��%  t�J& �t*$ �a� �7���Hc� & Hi�H  H���;f �q� �=�)  t����������%    �RHc� & �   ���%     �5�($ Hi�H  ��
&     �a &     �V���&     ǀ�;f     ���% ����v�   ������% ����   ���$Š[B �G($ ��   ��  �   �j&    H���% �SB ��D��W�% u1�*�E&    �($ ��uE�4�% �  H�e�% �SB �B   谾 �^��SB �R��% �   ��&    ���SB �5���% �   ��uH��% �SB �H��% TB ��
TB ��TB ��9  �=��%  t.H�=��% ��SB �A�����u�TB ��� ��yH���% TB X���&     ���% �����d�%    �USQ�=5^% 	um�-)�% H�:�) Hk�(H�H9�tH�   �(TB H���l�����u��]%    �xH�ߺ   �.TB H��(�F�����u���]%     ���TB 1���P  ��]% ����u:�3TB �-� ��~��&$    ��   �8TB �� �������m&$ ��   �   �=TB �T&$    �0U  ����   H�t& H��CTB H�\�H��������t.�ITB H���������t�MTB H���������u �   ��   H�H�����\B � ]% �O�VTB �x����CTB �oTB 1��g����ITB �oTB 1��V����MTB �oTB 1��E���ZH�޿tTB [1�]��O  X[]�S��TB �� ��TB ���� ��\% H���% �TB �у��uO��xH���%  PB �   �J%$ ��uH���% �TB �x��uH�|�% �TB �f��ubH�k�% �TB �U��x��xH�V�% �OB �@H�I�% �OB �3��uH�8�% �TB �"��uH�&�% UB ���uH��% +UB [�Ë�$$ ��\B H�0H��tH��9P�u�CUB 1��1����AU1��.0@ ATUSH���  ��M  �sUB �N  ��UB ������ ��UB �S  ��UB ���% �tS  ��UB �u�% �dS  ��UB �]�% �TS  �ǉ��% �� ��UB �=S  ��t
��%    ��UB �%S  ��t
��%    �=P�%  t
��UB �t���1��V  � VB ��R  ����   ��& ��   �Q�9�~+H��& H���  H�|��!���=�  Nظ
   ��
L؉޿VB 1������:*$ �d   �Ù���)*$ �'*$ �Ù���*$ �	*$ �Ù����)$ ��)$ �Ù����)$ �VB �����5� �4VB �����ZVB �nVB �T  �����T  1���@ �ZL  ��e �?   �����H�W�% H��u
�zVB �M  ��%     ��VB �L���H�-�% �WB 1�H���6���H����� 1��� �_����   �WB �XQ  ��tTH�1�H�hH��& L�,�Hk�A��H���\B  ��  H���\B I�} H���������u�Ic�Hk����\B �"$ �c�1Y% ��u�"$ 	   �L��u��!$    �;��!$ ��w��!$    �$��u��!$    ���u��t���!$    ��!$ ��w�=�!$ u��!$    �&��u!�=�!$ u��X% ����w
��X%    �>WB �� ��x�GWB ��������%    ��� �   �qWB ���% �P  ��u�   �{WB �P  ����   H���WB H�XH�A& H�<��{z  ��H�/& tH�4غ   H��$�   �x  �H�غ�WB �   1�H��$�   �P����WB 1�H��$�   �L���H��$�   ��� H��t���% �p�Hk�(H5�z) �H��& H�4�H�|$�	   �Ax  H��$�   ��WB 1�������   ��s@ �I  �3� �����=SW% �F���H���fS  �=s�%  H���% t\H�|$��[B �.   �= $  �u��WB 1��CJ  �=�$ u-H�\$H���   H���p� ��y��WB 1��J  H��H9�u߿�WB �M� ��x�I  �XB �A������XB �.� ��y�H�=��% �I  ��TB �� ��x��TB �� ��y��XB ������CI  ��YB ������K� �*N  ��E  �   �sF  � H  �  �   ��YB �i�%    �G�%    ���%    ���%     ��M  ��t$H�#& H�H�D�� �k�%    ��1��% �   ��YB �M  ��t.H��& H�H�D�� �0�%    �*�%    ��0���% �   ��YB ���%     �YM  ��tH��& H�H�|�������g�% ��YB �}M  ��t
�O�%    �   ��YB �M  ��tgH�]& Hc�H�=$ H�4�    H�<�u�����"�����0;$& �&�% }H�D1� ��0�k�% �
�_�%    �Y�%    �>RB ��L  ��~(���%    �3�%    �-�%    ��%    �   ��YB �eL  ��tH��& H�H�|���������% �
���% ������YB ������Zq  ��YB 1��������^ �ZB ������[ �3ZB ������J% �4�    ��J% �<�    蕱 �MZB �����W  �2����{ZB �����z<  ��ZB �r���蟬 �=�$ u��ZB �S� ��y
���%    �   ��ZB �K  ��t���A �   ��E  ��ZB � ����   ��ZB �VK  ��tH��& H�H�|��h,  ���%    �   �qWB �&K  ��t���%    H�|$�u.  ��   �{WB ��J  ��tH�|$�c0  �p����=S�% ��x'���  H��$�   �   H���s  H��$�   �'  �=�% t��Y�% ��% t�G�% �5��% �=��% �{(  ��]���듿�ZB ��\B �.���H��H�S�H��tH�s�WB 1�������H�� & �$WB H�4�1��E  ����1�9��^B u9��^B tH��H=�   u�1�ø   Ã�u'��u��u
�Ƀ������u��u	������ø�^B E1�98u,9pu'1���~0Mc�I��I���^B A9P|��~A9H����A��H��A��u�1��A��A��A�   �   D��D��D���m�����tA����A�A�ÍG����    F�1�9�`^B u9�d^B tH��H��Pu�1�ø   �1���w�   ��H��Q����ø�]B ��w
��H�� ^B �AVE1�AUI�������ATI��UH��S�=��%  ukA���9f  taC�<4 uZIk�R�P   ��_B � �e �q  Hc��% H��Hi�H  I�� ת% �=��%  Hǀ�<f  �e �����9f     t�..  I��I��u��=��%  H�-��% t����[]A\A]A^�(1  �   H��X��_B H��"H�D$�H  ��~�X4'    @�D$   ��_B �bH  ��~�84'    ��D$   �$ ��ZB �D$�#P% �D$�.H  1҅�~��_B �H  1҅���H�|$$�T$�E� ��TB �h� H�|$�����D$ �������_B ���% ��G  ��~
���%    H��X�H��x�=~�%  t
��%    ��`d �������% ��ZB �D$���% �D$���% �D$(���% �D$,���% �D$@�;$ �D$0���% �D$�[�% �D$ �Y�% �D$$�#�% �D$<�:G  1҅�~��_B �*G  1҅���1�H�|$�T$4������D$�T$���% �D$�?�% �T$ ���% �D$(���% �T$$�=�% �D$,���% �T$<���% �D$@���% �T$L���% �D$4�K�% ���% ��t
��_B �����D$H1�D���% �2`B ���% �5��% �����% 1҃����% 1҃��������% �6�% �����% 1��������% �T$H�q`B �p��1��������% ��~P�=��%  tG��u��YB ��E  ��`B ��u*�5��% 1���`B �N����=��% ~
�s   �k�����XB �1���H��x�U�   �A   SR���%     ���%    �-�%     ��K%     �iM% ����u�   �ϫ �WM% 1�D�2$ D�O�% D�<�% ��ad �   ��H�5��% H���% ���A��	u�8 u�@   E1���t
��A��DE�D9 u��uD9PuD9XuH�pH�H@�H�� H=�dd u�@��tH�5;�% H�,�% �>�%     �,�%     X[]�AVH�=�% �   AUATUS��� H���% E1�L��@  E��I������A���  I�H��H��@�   L���L9�u�A��@L��@  A�� 2  u¹�   �@  1�1��� ���% ��~|��
�   L�-��% A�
   �A�
   ��H�I�l L9�tRI��A�]���tF��
uA���6��A�^�:�����!��?w#H�H�� Bf �D��@  D��D��迬 A���[]A\A]A^Ë3$ �   �?   ��$ �������%     ���%     Hk�\���%    ���%     Hc��jd ���%     ���%     Hk�(H �d H���% �@���% 鏩 �{�% �ȉs�% ����  RH���% �z�t�B����   �h�%     �Z�% ���R�% H�H��H���`d  u
�8�%     Hc1�% H�����`d Hk�\���jd ��t1��� Hc�% ��%     H�����`d Hk�\Hc��jd Hk�(H �d H���% ��  H��0�d uFHc��% ���%     ���%     H�����`d Hk�\Hc��jd Hk�(H �d H���% �f  Hc����% Hk�(H�� �d H���% =�  �*  ��   =R  �   wA=�   �(  w=�   �  �   =�   ��   =   ��   �8   =P  �   =|  ��   w�k   =T  ��   �   =y  �   =  ��   ��   -�  ����   �   =i  wG=h  ��   =  ��   w�4   =�  ��   �   =�  �2=7  tg�3   =N  �=�  t[w�   =�  tR�   =�  tF�K=�  t8�3   =�  t1�6�7   �(�5   �!�   ��6   ��   ��   ��   1��� ��% ����   ���% Hc��% ���%    H���ɋ��`d tHk�\Hc�kd �Hk�\Hc�kd Hk�(�΃��5��% H �d H���% H= �d u=Hk�\��t	Hc�kd �Hc�kd Hk�(H �d H���% ��=�%  t<�������HcM�% H�����`d Hk�\Hc��jd Hk�(H �d H9?�% �T���H�2�% �@���t���% �
���%    X��V�=a$ u6�=��% 2v-1����;f  uHH  H=   u���=H�% ��   �������% �P���% ���% ��uY�����=$ ti��ueH���H�=}�% H���H��H��H�H�@H�   H9�v=�=��% �53$ �U�%     �S�%    u�   Z�w� ���%    �n���X�1��? u}�=#�%  t�   �Hc�% �
�%    ��%     ��%     H�����`d Hk�\Hc�kd ��kd Hk�(H�� �d H���% �R���% ��t�P1�荠 �   Z�Ã=��% u�m���1��ATI��UH��S1�M��tI��A�|$���u�ع   ������ہà   �>�B�����!��?v����H�H�� Bf � ��H���}���t6������!��?v
��H��u��H��߾�   H�� Bf D�"蘦 D���[]A\�S�   ��`B ��� 1�1�H���r� Hc��% H��H���`d �0���H���% �   ��@H��%�  H�g) Hk�HB�x�X=�Z& ��� ��   ��   H��t[�� [�� Hc�H�	�% Hc�HcD�H��<�t9Hi�@  D�F1�H�H�I9�tLi�@  D�TH��F����FH�t���AT�   ��`B USH����� �   ��`B H����� ��   1�1��@  H���C� ���% �   A�@  -�   ����    ��@  H�=@  DN�E1�A��?  D��H���
A������H��D��A������A��A��@  u΋n�% =i  ��   =�  w-�   ��`B �0� �D   �l   H���Ϥ ���%     �l-�  1Ҿ   �   ����F�9ԝ% }�   1��ߝ ���% ��`B �پ
   1�H�|$�ع���   H�|$�� �D   �l   H���W� H��[]A\Ë��% ��t��t
��uc�����t�����% ��u�s�����t ��t"��u;�=�$ ��SB �TB HE���aB ��aB P�   �3� 1�1�YH���ף ���L��% E1�1�L��% Hc�I9�t<C�C�<@8�t)v)�@��9�~�s�@��9�}C�<�C��   I��뿃��1�É�AW�   AVAUL�-��% ATA�ԙ��UH���% SLc�H���% L��M�H�D$�H���% H�D$�   A��A�����   1�E1�E��D9�~�B����y��B���   9���   �   ���Y�9�|��)�A��D�)��D��Mc�H�D$�1�M�LL$�E�Mc�M�M�H;D$�tfE�<AH��fE�8M����Hc�A��B��H�HD$�D��E�A��Mc�A)�1�M�M�L9�tfD�HH��fE�M���1�I����4���[]A\A]A^A_���1�H�5��% Hc�H�=k�% ��PH�=X�% �v� H�=d�% �j� H�=P�% �^� 1�Z�AUA��ATA��UH��SQ��   ��1ҍ	����� Ic�E1�1�L�A9�~0Ic�H�61�H�H�H�A9�~fD�zH��fD�L���H��E���Hc�H��H���H��X[]A\A]��� ��AT��U��H�=��% ��S��H�5��% �Hc��   H�=��% ���ډ�A���B���H�=��% ��D��1�A�   �)���1Ҿ   �<�    �� H�F�% �d  �   ���H�2�% �ډ�C9�~D�d  H��H�=�% �H�4�    A���D7�H�7�D���~�    �ƃ��t��������[1�]A\�P1Ҿ   � �  �� H��H�ؙ% �� 1�Z�ATA��1�U���   S��� �  H���L$�a� H��H���% �[� �L$D���L���% ���ĥ H��1�[]A\�AUE��ATE��U��S�V�=i�%  u*H��% D��D�Ɖ��N�%    H�/�% Hc����B 1�1���D��謞 �CD��D��H������B ��t��D��D�����%     Hc����B 1��=�%  Z��[]A\A]ËGGÉ�AW��   W�AVA�   AUATUSH��R���Hc��% H��HcҊ�
�9f �GHcX�$ �<� �e  u'Hc��$ �<���e  uHc��$ E1��<�D�e  A��Hc�$ A�   ���   %Hc��$ ���<� �e  uE1�<�D�e  A��Hc�$ �D�% �<� �e Hc��$ �4� �e ��	�	�u�e�%     ����% W�% IcŉN�% ���   E��t>1��t
Icŋ,��ed ��t
Ic�+,��ed ��~Icŋ��ed ��WtUIc�+,��ed �I��tHcЋ��ed f)S��tHcЋ��ed fS��~���ed 1�f)C��    t���ed fCHc�$ E1�<� �e  tIc�D�$��ed Hc��$ �<� �e  tIc�D+$��ed �=*�%  yIcŋ��ed A��tIc�D+$��ed Hc��$ �<� �e  u+Hc4�$ �<�D�e  uHc�$ �<���e  u	�=Η%  y
Ic�+,��ed Hck�$ �<� �e  u+Hc��$ �<�D�e  uHc��$ �<���e  u	�=��%  ~Icŋ��ed ��(  �CHc�$ �<� �e  u"Hc��% �<���e  uHc��% �<�D�e  t�KHc��$ �<� �e  u"Hco�$ �<�D�e  uHc*�$ �<���e  t�K��%     �=��%  ��   D�R�% 1�E����   Hc �% H��Hi�H  ��`<f H�;f ��
u�P|1�A��9� �B tH��H��	u�A�	   Lk�R�=;% D��$ D��Hi�H  A�	   A	����H���;f A�	1�H�H��	I��Hc�D9�tA�� �B ��u����P���wE��t̉�J�T: �<��;f  t���u���    t�~< t��C��$�B ���1�H�ŀ�B ��Hc	�<� �e  t�C����	ЈC�	H��H��u�Hc��$ �-�%     ����e ��tIcŋ��ed A�Hc��$ �<���e  tF+$��ed �=��$  �  ;��% ���% t:��~5���% ��t�x�% �=q�% u�K�a�%     �1�]�%     �%��% �O�% ��~�8�%     �2�%     Hc?�$ �   �<���e  uHcI�$ 1҃<�D�e  ��9��% ���% t:��~5��% ��t�Ք% �=Δ% u�K���%     �1���%     �%f�% ���% ��~���%     ���%     D%H�% ���% E��t�lE ���    f)S��u
���%     ��%     �n$ �T�%     ��D9�|	��D9�AL�9�|��9�L�  C�=M�%  t�A�%     �C��=~�%  t�r�%     �p�% ���Ȃ�C�=��%  t f�'�% fC���   0�)�f�Sf��% X[]A\A]A^A_�R��B ��, �=� $ ��)) u:�� $ ����w,���% ��B ��~����B ��B HM��- �R)) ��% �=$  ���% u
��$ �������%     �L<f 1����9f  ǀ�;f     t�z�u�B�   W�H��H��H  �����H��uŋM�% �=[�% 1ҋ5G�% ��  ���% �b�%     ���% �� � �e 1��   H�׺��e �=��%  ���%     �H�׹	   �@�e �   H���o�%     �i�%     �'�%     �m�%     �s�%     ���%     �o�%     �tHcP�% Hi�H  Hǀ�<f !�B XË��% ���% ��uW�? uR�5��$ 9wuG��u	�=a�%  u:���% ��% ����u1�Hcȃ<��9f  t���% �
9�uމ��% �   �USH��QA�% u4�=��%  u��u&���t�����  �{ �  �E  �9  ��t�=��% uC�1H���"  ���  H����~ ���
  H���!�����t���  H���o�������  �=��%  �t��u�C�S��1�)d�% �   ��u,HcC;)�% u�A�% �����(;�% u �-�%    ���t^����   ��uJ�2;��$ u���%    �f  =�   �[  �� �e    �K  HcC=�   �� �e     1��3  D�[�-f�$ 1�1�D�W�$ ���% A�   D����D��@�ǃ<���e  ��D��@ �t9�tA9�D�AD���ƃ��D����e H��H��u�@��t�V�% ���$ �
   �H�C��������% �C��������% �   D�SD���$ 1�1�D���$ �5	�% A�   D����D�����<�D�e  �� �tA9�tA9�D�AD���׃������D�e H��H��u�@��t�5��% �C�H�% �C�;�% �C�.�% �   Z[]�Hc�1��   Hi�H  H��<f H��H��0<f �   H���H���;f ���   ����Hǂ�<f     Hǂ�<f     �Hc�1��R   Hi�H  H���;f �L<f L���<f H��D���<f ��L<f H�      H���<f H��`<f �d�$ L���<f ���<f �U�$ D���<f ���<f �F�$ ǆ�;f     ���<f �4�$ ǆ<f d   ǆ\<f    ǆh<f    ǆ�<f 2   ���<f ��9���AULc�Ii�H  ATUSQH���;f H��u;1�9���  Hi�H  H���;f ���9Qu�V��9Qu1��~  H������nI��H�����������  ��tԋV�% ��~��H�<��6f 衷  �;�% �    ���Mi�H  ���I���;f Hc�H���6f ��% ����% �< �-   I��fA�D$��f��f������
��   tr��   th��   t`��ur�Z��   t6��   u^�=�K �5�+ �`��   t$��   u@�=Л �5�[ �B�=�[ �5�; �4�=�� �5�K �&H�}'% Hc��<��4���B ��7�B 1��)$  1�1�I�E k��'   k�����a�  Hc��% Hi�H  ���;f t�#   H���� �   Z[]A\A]�H���������AUATUS��RH�5��% H��_f H��H��A����Y�B 1��#  A�   ��T  �ߙA��Hc�Hk�
H�ŀ_f H���������t��H��f�]�A��u�Hc�Hk�
H�� `f X[]A\A]���  �=��%  u�/�%    �AVAUATUHc�Hi�H  �=��%  SH���;f Hǀ�       t[]A\A]A^�!���Hk�
��E1�H�� `f H���0�����uNMk�
��I�� `f L��������t,Ic���L��A��Hk�
f��`f �W�  [fD��`f ]A\A]A^�I��I��u�[H��]A\A]A^�-�  �p�% 	   ��5�%     �[�%    Ã=�# u"P�~�B 藹 �<�%    ������% Z��%�%    �   ���% �QE1���%     B�<��9f  tD���/���I��I��u�=-%  t�e����=��# Hc��% ��t-�=��# 	u��u���t��	t"���u���%    XÃ�t2��t-��	u(�q�%    ���%    ���%    �+�%    Hc��% �5.�% I��Hi�H  �� =f �4�% Hc�% �J�� �% �H���% ��uC��t)��t����   ��%    �   ���%    �w�p���   G��5��% �a��t���%    �Q��	uF��t)��u@���%    �4��t��u*���%    ����%    ����%    ��z�% ���%     �5��% �5h�% �5��% �5`�% �52�% �5X�% ��uHc�k��dd #���Hk�
H�k� ed #�k��dd #D�-�% �53 & ��;f 1ɉ�% � Af �<��9f BlH���p8H��H  H��(�8�z�@�x�z��x�z��xH��u����%    � Af �:�%     ��*%     ��n � Af Z鑲 ���%    �\�% ��tHc	�% Hi�H  ǀ =f    �=%�# u*�1�% ��w�   H��@@u� � �t	��t�i����P�)�% �#�%     �����% �������%     ���%    Z�PH���   � 8f �L  ���%    Z�P�    �=ņ% � �e �bL  ���%    Z�ATUS1���  �=��% H���E�  ���B H��I������H���% H��u6���B �!O  ���B H��H������H���% H��uH��H��B �c  �j�%     � �e �c�  �3�  ��  ��  ��  ��  �=��#  t H�=/�% �b���H= � ~�ʀB 1��  H�=�% �¡��H��tH��H���B 1���  L������L��H�������    �|�B � �e ���%     �AK  Hc3�% []A\Hi�H  Hǀ�<f D�B �G* �=�% �5��% ���% �t�%    �AUATA��U��S��Q�=��%  t���%     �p� A��A�   EN�=��# v��t�	��~)�����"�   ��   �=��#  �   D���   ��~��	~�=��# �	   E���   �tN  �   A��1��=��%  ���=��%  ���% u�v�% A��~9��tk1�Ѹ��d H��(H=  u��)$    ��	$    �y	$    �7��u21�Ѡ��d H��(H=  u���$    ��	$   
 �@	$   
 �=��# ��% ���%    ��%    �M�%    ���%    ���%    �{�%     �y�%     �'%     �U�%    �-��% D�-��% u��B ��~(����B ��B HM������B ��wH�<ݰ�B � ��) X[]A\A]�/���S�P�B � 8f �d�%     �Ǡ��H�h�% H����   �]�%     �4�  ��uH�=E�% [��������% �5��% �=��% �/�% �����$�% ��  �I�  �?�  �0�  ���  ��u
�S�B ��  H�=��% 衞���=vl&  t�/ [�|' [�P�4�% �5�% �=@�% �:�%     ���%     �:�%     �`�%     ���%     H���%     �]�%     �K�%     ���%     ���%     ������<�%     Z�U1�H���H��SR1����%     �H��H��H�^�   ����� H��H�麅WB H��H���% 1��   ��J  �   �`�B �w  ��tH���% H�H�|�������
Hc؉�1Ҿ   蝵 �%�%    H�H���% H���% X[]ËB�# �j   ��t.��t�k   ��t 1�������l�P�i�B 1��`  �j   Z��R��_B �.  1҅��-�% ���҉m�% H�>�% H�'�% tH�BH��% �o��x���H�	�% H�JH���% �H���% H�PH���% ���% �H���% H�PH���% ���% �H���% H�PH���% �x�% �H���% H�PH���% �f�% �H���% H�PH���% �h�% �H�s�% H�PH�h�% �F�% �H�Y�% H�PH�N�% �l�% �H�?�% H�PH�4�% ���% �1�H�#�% ���9f H��H�rH�5�% �
H��u�X�H�=}�% ���%    �AT�   H�=d�% US���%     �� H�PH���% H���% ��!���9�u���%     �o��ou���%    �^�C���w
H�,���B �4���B ��v*�عd   �   ���e ����e ��A�Љ����B 1��(H  ����H��޿��B ��1�芛��H�3�% H�PH�(�% H�P�H��% H�P�hH��% H�PD�`H���% �P���% H�PH���% �P�Ȼ% H�PH���% �P���% H�PH���% �P�ֺ% H�PH���% �@��% 1�H���% H�JH���% ����9f H��H��uۃ=��%  t��%    �A�%    ���_B �-  ��ܿ��B �  ���D�������#     �������#    �Z  []���%     �4�% A\���%    �SH�����B ��  H�b�% [�k�% �u�%    ��+%    ���%    �Q�=X�%  tK��  �5��% +��% ���B �6�%     �*ȉ°��%     �*��Y� �^��Z��f  �=��%  ��   H�=��% �� �=O�%  ���%     ��%     ���%     ���%     �Y�%     H�R�%     ��%     �ڹ%     ��%     �b�%     t��  ������   �g�?�% ��t]H���% H�PH���% � �H�5��% H���% H�=y�% H)��?  H�=��% ��� H�5^�% 1��ÂB ���%     �g  1�Z�H�]�% �8�u����H�PH�H�% ��H�PH�9�% �P�WH�P�=�%  H�!�% t"�PH�Hf�WH��% �@��	�f�W��@��f�GH���% H�PH���% � �G�Hc+�$ AVAU�<� �e  ATI��USt�����H���% A�$H�HH���% �H���% A�L$H�rH�5��% �
�=m�%  H�z�% fA�L$tH�rH�5g�% �
fA�L$H�W�% �f��H�rH�5F�% �
A�L$H�8�% �
H�W�% H�(�% H�Q�H9�vy�=x�#  t[]A\A]A^�M���H��H+�% 1Ҿ   D�4D��Mc��Ϯ L�-��% H�5��% Hc�H��H��I�I)��H�=��% ��� H�-��% L�L�-��% H�-��% [L��]A\A]A^�2���AUATUS1�AP�<��9f  tHi�H  ���;f u���!���H��H��u֋T�% �B���ts��w��$�`�B ��������r������������`������6������ �����>���������믿ԂB ��� Hc��% ���%     Hi�H  Hǀ�<f ��B 뀋�% ��   ��;f 1ۙ�=�% ���Lc�<��9f  �5  H��L�mH��H˾% �=(�%   EtL���'����=��%  tL�������}2~���;f    �s�% �u[���   ���9�uL�<��;f  tBH��`jd ��B �P   1����e ��A  Hc��% ���;f     Hi�H  Hǀ�<f ��e �=��%  t{�=��%  ur���% �ș�=��% ��u_���   ~%H���uH��B�� �9f @8�t���B 1��  H�E H��tH�ڋ@H��B��"�9f �H�؋T�% H��B�� �9f H��H��H  H�������1ۃ<��9f  t{Hi�H  ���;f ��yj��<t<t%�]���% ���ȉ��% t�y �A�<y �:�=�w%  u�    ��B � �e �=  ���;f ��%    ������w% H��H���n����=ſ% u�=��% t��� ���% ���% ��t5��t��t8��u?Z[]A\A]�-������  �*n 薢��_[]A\A]�  ^[]A\A]魠 Y[]A\A]����X[]A\A]�ø   �G H�� H�Ghø   �7H�� �WH�OD�G�G H�Gh�HcWh1���Pt�B�GhH�@�t�D �   �Gl   ËWh1���t�ʸ   �WhHc��D �Gl   �AVAUE1�ATA��US�/H��D9kh~YB�|+����< t:�ЋK<_w09�,)�H�CHc�H��D�2A�A��@  �s��D���T~ �����?  I���E��t0�_   H�S+CH�H����=@  �s��[]A\A]A^�~ []A\A]A^�AUATUSH��R�=;%  t�Cl����   �ȉCl�~�= \&  t�l t�H�G�oH� Di�@  D�hA�ŋCD�9�~���A& 9�
�A& 9�
�@  D����5�[& D���� �5�[& B�<&=�^& � ��A��@  �X[]A\A]�H�D$���  E1�Ǉ�     H���  Ǉ�      A9�}=I� A��H��p�@�w�L�G���D�O�A���G� A���G�    �G�   A)�D�_��Ë��  ���  �����  9�u
Ǉ�      Hc��  Hk�pH��@h    �@ �@l   1�9�~Hk�pH���Dl   ���I��I��I������H��t!A�2@��tIc��  I��Hk�pL��`�����A�1@��tIc��  I��Hk�pL��?������H���  �8 u�UH��S1�R���  9�~!���  )�y�Hc�1���Hk�pH��K�����X[]�U1�SH��R9��  ~2���   tH���  �8 uHk�p�Dl   Hk�pH��H�������H���  � ���  X[]ø   L�OxH�� �7Ǉ�      �WH�OD�G�G H�Gh�Gp    ËGp9Ght�����H���Ah9Apt
H���x�����ø   �G H�� �Gp    H�Gh�H��I��A�0@��tH��I��������Ah�Ap�SH��@���[����P���?w��H��������<uH���r����   �<����[�H�Gx�8 t
�   �
����S���    H��tH�Gx�8 u�Gl   H������H�Cx� ���   [�S1�H���K!�ĄB �	   1�H�|$�ҍ���   H�|$貣 H�� Bf H��H��?u�H��[��Bx%     �USW�=7x%  t
�+x%     Hcķ% RA�!   1�h�e A� Bf �   1�Hi�H  �@�e ��y%     ���%     ��y%     ���%     H�;f H�}% �b���H���% ��   1�� Bf A�!   � �e �@)��r�����% Y^��t(��tB��t=��t��t>�΄B ��uG�R�% ���2�S�% �ȍ�<�% ��H�H���hd ��(�% ���	��% ��?H�H���ed �=��# 	u��% ��H�H���hd �3@��t� �e H���������H���% A�Bf A�!   1�� Bf �`�e � �e �@�e �P������H��A�D�e E1�1�1�1�H�È   �����H9�u���v%    X[]�Q�@�e �B����`�e �����=�%  t1�� �e Z����X�P�@�e �Y����`�e ����� �e Z�9����Cv% AVAUATUS��t�ȉ/v% u�x%     �x%     ���% ����$ thH�N{% H���   H��tU�=�w%  t��tH1��@�e �>���H�"{% ��w%    ��u% �   Hǀ�       ���% ���%     ��w% �=V�%  ��   1ۃ<��9f  ��   9�% ��   Li�H  E���;f E����   A��D��@�e �   Hi�   A��L�� �e L����������   A��uz����e  ti���% ��@�e ��9�t��uQH�4�`jd H��4�e �@�e �N����=��# �l   ��v%    ��v%    ��t% �   t�W   1���m L���U���Aƅ�;f  H��H������[]A\A]A^�Hc�s% �B��;�s% uH��y% Hǀ�   ܄B �@����e ��s% Ë�s% 1�9�s% tHc�������e ��s% �USQ�G=�   �}  �=�   u1������as% �b  ���Z  �=پ%  �T  ;i�$ u��u%    ��s% �   �6�=��%  �"  �w;5+�$ u(���%    �`�e �Q����   �����   ��  ��% �% �% �% ����   �=
�% ��r% 1�1�H��x% ;4�@Df ��   �<��9f  t.9�t.��t��r% ��%    �`�e ������{@���t���9�uW����Hǁ�   �B �A��Hǁ�   �B �/��Hǁ�   �B ���Hǁ�   $�B �Hǁ�   6�B �H��H���S�����t��q% 1���   �=�q%  tk��0<	w��ȿ   H�4̀jd ������>@��tH����   ������Q   � �e �/�%     H�4̀jd ��1  H��w% Hǀ�    �e �����o�`�e @��������Å�t	@���|���@��u;�=�v%  �Լ%     t8�Q   �t�e � �e �1  H�#w% Hǀ�    �e �@��u
���%     ��Z[]�����U���e �v�B ��7e S1�H��(�;  ��7e ���B �,  ���e ���B �  ��7e ���B �  ��7e ���B ��
  ���e �ǓB ��
  �|�e �ٓB ��
  �x�e ��B ��
  �ٺ�B �    H��1����4  H��H��H���
  ��
u�H��([]�AT��B US��  �&�B A����  �-�B ����  E��H�=š%  u?�Ņ�5�o�$ ��t��u������H�v%     ��H��u%     ���~�[]A\�H��u% H��tQ�PH��u% H��tH�@Z�X�H��u% H��tH�@���H��u% H��t�` 1��H��u% H��tQ�P(H��u% H��tH�@`H��tZ�X�H�pu% H��tH�@`H��t���H�`u% H��t(���   ��   Oу��   O�1Ʌ�Hх�H��`0�H�+u% H��t/���   A��   AOȃ�A�   AO�E1���AHȅ�AH��`81��H��t% H��t�`@�H��t% H��t�`H1��H��t% H��tH�@PH��t�����H��t% H��t�` �H��t% H��t�`(�H��t% H��t�`0�H�yt% H��t�`81��H�gt% H��t�`@�H�Wt% H��t�`H�H�Gt% H��t�`P�H�7t% H��t�`X1���UH���   S��P�)���H�2t% H�(�XH�PH�!t% Z[]��AT1�H���E1�U�#   SH���H��H��H��H��)�A9�}�    A���������H��[]A\鷅��S�K   �=   �ׄ����u�
   [�Ȅ��H��H�|$�����H�|$����������6�B �q���H���1��SH��s% H��t�H�[��[�AUATUH��SH���  H��$(  H��$0  H��$8  L��$@  L��$H  ��t@)�$P  )�$`  )�$p  )�$�  )�$�  )�$�  )�$�  )�$�  �=�r%  tH�5
% �L�B �K����
��r%    H��$   H�=�	% H�T$H��H�D$H��$   L�d$ �D$   �D$0   H�D$����H�5�	% �z�B ����H�=�	% �o�����   L��H��H��$   �   �D$   H�D$H��$   H�D$1��H�L$L���D$0   �[/  H�-r% H��t�} t�U H�m��}�B �s  ����   ���B ��������   L��H����H��H��H�|輁��� "H��L�hA�$��t&�󿫕B �]���H��tA�E \I��A�] I��I����fA�E " ��H��H����H��H��H��!H���`���I�蹰�B H��I�ĺ��B H��1��.  L���k���L������H��������AT�   UH���ՕB S�   �C  ��~H���% H�H�|��ׂ���É����} Hc�����I��H��u�s��ٕB 1��m����U H�ƿ�B 1�謁��L��[]A\�AWAVA��AUATUH��S��H���=�$  ��   �   �+�B �ի$     �  A�ą���   H�H��% �3�B H��L�<�L�,�    L���x�����uH���$ h�B �:�B L���\�����uH�}�$ X�B �o�@�B L���>�����uH�_�$ H�B �QI��E1�A��D9%l�% ~3H�k�% I��J�<(�?-tH�t$I���E(  �D$A����e I��
u�H��$ ��e A��tA��t51�A��ugH��$ ��E �SH��$ �C������	�f�E �4H�Ī$ �C�K��
����	ȉ��
	ȍK�
��	ЉE �   H��[]A\A]A^A_�1��� Q1��� �=%o%  u�o% +o% ��  1�k�#��Z�Q1��� �=�n%  u��n% +�n% Z�鮢 ��AVI��AUL�-E�% ATU�-4�% S�   )�A��9�~I�t� L��H���ŀ����u��E1�[D��]A\A]A^�1��P�����Z��������H��% S�/   H�H���~��H��tH�XH��[ø����H��H�H����   �H�G�9w~�w�9w}�w9W~�W�9}��H���1�H��D�G(�H��H��E��~	H9J v1��H�B0H9�s1�@84uH�HH�J0�B8    ��B8A9�~-Hc���@�t
<�B81�H���H���H��H��H��H9B0r�D;B8��B8    �   H�B0    �H��HcO(H�w<H����AVI��AUATI��U1�SD�oA9�~H��L��H��H��I$H�3�&}����u��1�H��[]A\A]A^�UH��H��� Ge SQ����H��H��u$H�� 8e ����H��H��uH��r�B 1�����H��Z[]�H���?0u�xuH��H�T$��B �
H�T$���B 1��||���D$H���H�=�l% H�5�l% ���Q�   ���B ������t#H���% H����B H�t�1�H�5�$ �M}���H�5|l% H�=ݳ% 1�1��Q(  H�Ͷ$ H�5ƶ$ ���B 1��}���   �ǖB �P�����t"H���% H��ԖB H�t�1�H�5��$ Z��|��H�5l% H�=w�% 1�1���'  H�g�$ X�SH������H�X�@   [�UH��SQ����H��1�H��t|�C��tu�{�   wj�C�$ŀ�B H�[H����{��H��JH�[H��������:H������1҉C��w	H�����B H�C�S��H����|��H�C�Z���   Z[]�Q����1�H��t�x t�xwH�@���Z�Q�����1�H��t�x t�xuH�@H�H��Z�R����W�H��t�x t�xuH�@� X�RH��t	H�=A�% ��   �z��f� . H�)�% H�5"�% �> t���B 1��q{��H�=
�% X�!  H�=��% �? u
�|�B ��z��S1Ҿ �B 1��\&  H��H���b!  H�޿*�B 1��%{��H��[�P�XRe �y�B �K����TRe ���B �<����PRe ���B �-����LRe ���B �����HRe ���B �����DRe ���B � ����@Re �ԟB ������<Re �ݟB ������8Re ��B ������4Re ��B ��������e ��B ������Qe ��B ������Qe ��B �������e �9�B ������Pe �C�B �y�����Pe �O�B �j�����Pe �X�B �[�����Pe ���B �L�����Pe ���B �=�����Pe ���B �.�����Qe �ޙB ������Qe ��B ������Qe ��B ������Qe ��B �������Pe �B�B �������Qe �M�B �������Qe ���B Z�����P�0Re �ҞB �����,Re �ܞB �����(Re ��B �����$Re ���B ����� Re ��B �x����Re ��B �i����Re �c�B �Z����Re �o�B �K����Re ���B Z�;���P�Re �ɞB �+�����Qe �-�B ������Pe �c�B �����Re ���B ������Re ��B ������ Re ��B �������Qe �&�B �������Qe �;�B �������Qe �M�B ������Qe �d�B ������Qe �q�B Z����P�Re �ɞB �T�$ /   ���$ a   �ļ$ �   ���$ �   ���$ �   ���$ �   �H����$Re ���B �9���� Re �ǟB �*����Re �|�B �����Re ���B ������Qe ���B �������Qe ��B �������Qe �*�B �������Qe �6�B �������Qe �A�B �������Qe �L�B ������Qe �X�B ������Qe ���B ������Qe ���B ������Qe �-�B �v�����Pe �c�B Z�f���P��Qe �x�B �V�����Qe ���B �G�����Qe ���B �8�����Qe ���B �)����|Qe ���B �����xQe ���B �����tQe ���B ������pQe �̜B ��������e �؜B ��������e ��B �������Pe ���B �������Pe �ΙB ������Qe ��B ������Qe �0�B Z����P�lQe �؛B �����hQe ��B �s����dQe ���B �d����`Qe ��B �U����\Qe ��B �F����XQe ��B �7����TQe �ɛB �(����PQe �-�B �����LQe �=�B �
����HQe �L�B ������DQe �Y�B ������@Qe �f�B Z�����P�<Qe �W�B ������8Qe �i�B �����4Qe �u�B �����0Qe ���B �����,Qe ���B �����(Qe ���B �����$Qe ���B �r���� Qe ���B �c����Qe �КB �T����Qe �ߚB �E����Qe ��B �6����Qe ���B �'����Qe �	�B �����Qe ��B �	����Qe �)�B ������ Qe �8�B �������Pe �I�B �������Pe �[�B �������Pe �j�B ������Pe �x�B ������Pe ���B ������Pe ���B �������e ���B ������Qe ���B �s�����Qe ���B Z�c���U��Qe �����B S1�H��(�J���H9�t,�K���B �    H��1��y   H�4�@Df H��H��������H��([]��Hc�Hc�H��H��H��É���������1�)Љ�1���)�9�|��1�������Hc�Hc�H��H�H��ø   +��$ ���$ Hc��% uHi�H  Hǀ�<f ֣B �Hi�H  Hǀ�<f �B ���%    �P�   ��B ��%    �� 1�1�YH���^ P�   ���B �� �   �^   YH���}^ P�   ���B �ć �   �`   H���[^ �   ��B 裇 �&   �6   YH���9^ P�   ��B 耇 �&   �6   YH���^ H��  ���  H��   H���  H���
����ԩ%     H��  �USR�   �=��% Hc����%    Hk��0Ef H��`Ef H���\  ��B H���q����uƃ`Ef  1�H��H����H��H��H�ȉs�% X[]�USR�F�# �Ȩ%    ��	wK�   H��@  uY��  uc�>t1��   ��   �J  �=�# Eظ  ��B E�TB HE��=�$�B 1���   �J  �%�����SB � ��   �J  ��B ���   �J  ��B �   �$� 1�1�H����\ f�-��$ f�}�$ X[]Ë�$ ��t��t
���t����������$ ���$ �<�    ��V ���$ ��t��t
���t����������$ ���$ �<�    �sV R�=ƽ$ �   +5�_% �5�_% � �=�_%  Hc��% uHi�H  Hǀ�<f ;�B �Hi�H  Hǀ�<f G�B XËr�$ ��t��t�1�Ƨ% ��~'���ʉT�$ ����% �����=�$ ���% �5q_% �=+�$ �~  ��t��tË�$ ��t�����$ ������$ �9=q�$ uE�=(�%  u=R���% �����=&�# H�u	�4�`Re ��4��Re 1��R �i   �����X���,���9=�$ uP�=�% ������   1�Z�LR �9=��$ u%P�?�% �   �   �p�i������%     Z��9=β$ u!H�Ŧ% f���% ���%     f�P$�9����ATU�`Ef S1�H��   ���@�  �   H��H���(  �P�B H����o��I��H��u$�   ��B H���  H��H��fǀ�Se   �-H���   �   H���o��L���n��H��H��fǀ�Se  H��H��H���r���H��   []A\�ATU���   S���R�B ��D���   �,� �{���H����Y �   �[�B �� �߉��H���Y D9�uݾ   �d�B �� ���[H��]A\�Y Hc�SH��Hk���H��`Ef �����=f�% ��H�%     u�T�% [�9=T�$ uP�=C�% �����   1�Z�P �AWAVA��AUE1�ATA���   U��S���m�B AP�_� ��D���H��A����X A9�}&�   �v�B A���5� D��D��A��H����X �Յ�    �   ��B H��� D��,�H���X �   ���B �� B�<�D��H��X[]A\A]A^A_�xX P�   ���B 迁 �&   �<   H���VX ���$ �   �5�$ �=�$ ���������$ �   �5ͳ$ �=ĳ$ AX��0�����P�   ���B �Y� �   �l   H����W Hc�[% �   H�<��B �.� �5��$ �=�$ H�� �ǯ   �W HcA�$ �   H�<�ЧB ��� �5´$ �=��$ H����x�W ��$ �
   �5��$ �=��$ ��`�2����L�% �	   �5z�$ �=q�$ AX��@����UH�����B S��   P���|� �U"�} Y�t���
[H��]�W UH�����B S��   P���H� �U"�} Y�t���
[H��]��V ���% H�=�% � �%    �&�% H�5��% �	�% ���%    Ã=c�%  t1�1����B �HHc��% ��y1�1���B �2Hk�P��B �P   ��Df 1�H��`Ef �i���   ���@ Y��Df �j����=&�%  u�"   1��}M �=�%  t1�1��Z�B ��   �L�@ ���B �-����@_d P� _d �   ���$ �����`Ff HEȋ�% �����   1�Hc�H�Ѻ��B �(i���   ���@ Y�`Ff �������u�   ��@ �եB ����P�ߠ% �   �p�����`�%     Z��Ƞ%     �Π% �H�% �ATH���1�U1�SH���H��H��L�d�L9�t)�;�j����!��>v���H�H�� Bf � �H���҉�[]A\�H��% H���I���p1���H��H��H��1�H��H9�tA�<
u�H�����AVA��AUA��ATI��U��SI��A�|$���tE��
u��D��A������i��A�^��!��>w�H�H�� Bf �D��@  ��D���mT ��[]A\A]A^�U�   ��B �`Ef S1�R�} �   �H   H���7T �5ڮ$ �=Ѯ$ ��,����5Ů$ �=��$ H��H��ރ��3�����`u�X[]�U�%�B �`Ef S1�V�   �8} �   �H   H����S �5r�$ �=i�$ �������5]�$ �=T�$ H��H��ރ��������`uǃ=��%  t<Hc=^�% H��Hk���H��`Ef �����5�$ �-�B �=�$ Y��[]����X[]Ã=2�%  u"�&�%    �@�$ H�1�%  Ye f��% �AVAUATUSH��P�=n�%  �h�%     ��   H�=/�% 1�H���������   ����؃�df��V% H�	�% Hc�Hր> ��  1�H��H��E1��H��H��H��E��I9�s0A�,�<

I��u�P   H���9  A��OwB�, A�n�)A����I��P   L���  1�H��L���H��H�Ѝl�H��������   �5V% ���H����f� ��f��U% �Q���H�"�% f�@f�U% �2����=�%  ��   H���% H�PH��t1���H��% 1ۋP �(f��U% f�P"f��U% 9�vIH�ŝ% H��H��Hx� t$H���   ��z �5iU% �=`U% H���Q f�RU% H���H�Y�% �   H�<� Ze �z H�b�% �7�% �=U% �R"���� �t
�H���6Q H��P[]A\A]A^���%     ËG$H�=�% f��% Ã=͏%  t1�1��/�B ����P��Se �����Z�B����=ɘ%  u1�1��d�B ������=ސ%  uP��Re ����Z����Ã=��%  u�"   1���G �=��%  ubQHc��% ��y �6����������Re �V����j�% ����Z�Hk����B �P   1���Df H��`Ef �c���   �Ɵ@ X��Df �[���Ã=�G%  ATUH��S�t-��t��t1���  �G;*�$ t;ڧ$ u������  ��uS�=қ%  t2�==�%  t)H�=�% ��@ u�=Ч$ �T����w  9��$ �H  1��   ��F 1������S  ����   �����;nS% ��   �} ���$ x�����t���$ ��������AS% �} y�e�$ �t�W�$ �������S% �Et�5�$ �������S% �Et��$ �v�������R% ���$ 1����e  �}�����W  ��$ �D�������R% �*  �} �$  �'���;�R% �  ��R% ��R% E�J�wR% 9�}���$ ��������cR% �UR% ���'�����9�~)���$ ��������:R% �,R% ���#R% �!R% �R% �R% E�J�R% 9�}�7�$ ��������Q% ��Q% ���$��9�~)��$ �`�������Q% ��Q% ����Q% ��Q% �Et�֥$ �1�������Q% �}��t(���$ ��������Q% 1���}  �|����]�}����m����=��%  �  ��t@��t����   �`�S�% ���  Hc$�% �ȉ<�% H�Hk�Ƅ`Ef  ��  Hc=�% �   �0Ef �F�%     Hk�H��`Ef �
  �  HcҘ% � �%     H��Hk���`Ef  ��  �Q����  �={�$  E��b��A�č@���?�m  Hc-��% ���]  Hcu�% Hk�H��`Ef H���/���=�   �8  �ED�$+�j�% H�� �   �=��%  tV�=��%  t�� t��t9M�$ t9A�$ �!������%     ���% ��% H�b�% H���  ������  �=I�%  t9��$ t��t9�O% u
茹���  �=Ɨ%  ��  9��$ u��$ ��% �����1��9��$ u!���$ ��% ������   �����Q  9��$ u#�3����`Ue ��Ue �=K�# HE�H�l�% �b9X�$ u����1��   �B 1��^�����  9/�$ u�����1��   �uB 1�������  9�$ u����H��% �Te f�ۖ%   �2  9ܢ$ u1������  9Ģ$ u�   1��B �����y  9��$ u1��   ��A 1��d����Y  9~�$ u1�������  9f�$ ������   1���A ������#  9<�$ uV�dy% �    �   ��RB ����O�Hc�% �@y% H�Hi�H  Hk�H Ze H���<f �ps H���7 ��  9*�$ ����������6  9�$ uQH��% �5ĕ% 1�� ��9�}�V1��   f���% �A H���% H���% H��HBf�8�t��V  9��$ uOf�r�% �B�f��uH���% � ��1��   f�Q�% �@ H�D�% H�a�% H��HBf�8�t���  9X�$ uSH��% H�7�% H��HBH�x ��  f�8��  1��   �W@ H��% H���% 1�H��HB�\9��$ u\H���% H�ܔ% H��HBH�x �z  f�8�p  1��   ��? H���% �   H���% H��HB�P�@  9��$ uYH�[�% H�x�% H��H��HAH�PH���  � f���  f�y$f��u�   �Ҿ   ��   �Ҿ   ��   9D�$ u&H��% f���% f�P$��%     �   �   9�$ u7H��% f�Ɠ% f�P$H�@H����   H�ғ% �@$f���% �   �k��u���   t���   t���   ��������5s�% H���% �FD�Hc�H��A9�~L�IE�LH�� A9�t����1��4f�7�% �   1��> �   �#H��L�@H��HQ�R9�t�L��9�}�����[]A\ÿ�Te ������=υ%  t�=��%  u1�1��ͦB �����=ì# t�=��# 	�@Xe u�`We ����R���# ��u��t1��B 1�1��������Ue �'��~��uH�5a�$ �k�B �[��1��=ۑ% �`We X�^���� Ve �T�����Ue �J���� Ye �@����=/�# w�=*�# �`Ue u� Ye ����f�F�% ��f�=�% f��f�5�% f�'�%  ����%     ��$ H��%  Ye f�ؑ% �z�$ f�ˑ%   f��% 
 ���=��# ���% �"�%     H��%     ��%     ���% ����u6f���$ ([�$ f���$ (\�$ H�ɣ$  Ye )�$ )#�$ �=<�# wf���$ þ�  �HZ��Q�w�B ��Z��H��tH��� Y���   �dH�%    H��# �<  ����Z�ATUSH���nY���   1�H��I���Z��H���TY��L��H��1�H���Z��H��[]A\�ATI�����B U��S�IZ��H��1�H��t&L��Hc�H�پ   �,Y��H��I���X��1�D9���[]A\�AWAVI���P�B AUATI��USQ��Y��H��H��uL���B 1�����H���@���1Ҿ   ��H���Op Hc�H��   H��I���Y��H��I���X��D9�~L���B 1��3���M�.��Z[]A\A]A^A_�UH��1�H��S��B H��Q�;W����u�   �F1�H���B H���W����t�1�H���B H���W����t�1�H����B H����V��������Z[]�ATH���1�H��UI��S�H��H��H�\2�H9�uI�$    1���{�/t�H�����X��A�,H���<+@��t"@��.tH��u�L��H�޿�B [1�]A\�W��[]A\�SH���;@��t�`X��H�ÈC���[�AWH���1�AVAUI��ATE1�USQH���H��H��H�,H���H��H��H�9�r-I��)�E1���E��H��L��M�L��� W����tA��D9�s�E1�ZL��[]A\A]A^A_�USH��Q�wV��H��H��uH��H���1��E�B H��H��H�r�����H��Z[]�H��t6H��SH�R�H���D� ��V��H���I��1�L���H��H�Ѐ|� [�����1��AW1�E1�AVI��AUI���ATL��UH��H��SH��H�$H���H��H��N�$)L���H��H��L��H����U��H��tH�<$J� L��D���H��H��L)�H���H���$U��I��I��H��uR�m�B 1������_L��L��H��L$�U���L$��u3H�4$L��H��L�����H�<$1�H����H��H��I�H)ˊM ��u��A�H��I��H����A� H��L��[]A\A]A^A_�H���1�I���H��H�y�H9�HG�H)�L�����H���1�I��H���H��H��L�H���H��H��H�I9�vPL���bT��Z�������1��I���1�I��L���H��H��J�	L���H��L�H9�rPH)�I�<��S��Z�������1��AT1�I��USH��PH�L$8L�D$@I���H�t$(L��H�T$0L�L$H�H�D$p�D$   H�D$H�D$ H�D$1�H��H�Ӌt$��/w��H�|$ ��H��t$�H�T$H�JH�L$H�:H��tL���H��H�\��H���WS��H��H��u���B 1�������fH��L��H���Z���H�D$p�D$   H�D$H�D$ H�D$�T$��/w�Ѓ�HD$�T$�H�D$H�PH�T$H�0H��tH��H���C�����H��PH��[]A\�H��1ɾ(�B �ɨB 1������1�H��t'UH��SH��AP�3T����xHc�H9�w�D� �C�Z[]��H���   H�L$8L�D$@L�L$H��t7)D$P)L$`)T$p)�$�   )�$�   )�$�   )�$�   )�$�   H��$�   H�L$�D$   H�D$H�D$ �D$0   H�D$�O���H���   Ë^B% �����SB% ���B ËIB% �����>B% ���B ��(B%     �"B%     �1�H�<� Gf  uH�H�<� Gf �H��H��u��S1�Hc�H9<� Gf uH�G H�@h    �"�  H�� Gf     �	H��H��u�[�USH��QD�O8A�����   A���&  �W,�w0A�   1�H� �(  ���ϭ% u�{tAH�C �   H�x0��4 ����   �C��w��s4��t
��   ���ZH��[]�?�������   H�C �   H�x0�4 �C8�����   �O4�W(A�   �w0H� �'  ���>�% u�{t'H�C �   H�x0�=4 ��u7�{wP�C�$��B ��u"H�C �   H�x0�4 �C0   �C8   ���u�K��w�   H��,t�C0    X[]�1�H�� Gf H��t�O9H<u�x8 u�H@H�@C�@ �H8H��H��u�ÍF�AWAVI��AUATA��USQ��w����I�      1�A���D��L���P�  A�Ņ���   Ic�H��H-M�% H�}h u�1Ҿ   �H   ��g H��H�����  H�]hH�CC�@ H�k �C4    A��wiD���$��B �E�C,�E L�{0   �C8�����C(�A�E�C4   �C,�E E���C8������   EC(�H���j�  �C8   �C,�C0   �ED�cH�߉C<�   ��������Z��[]A\A]A^A_�1�1�H�� Gf H��t'�w9r<u�r8��t�r@�   H�B    �B8    H��H��u��D�O0E��t*SH��A�����   �  A���(  A��th�{  �O8�t  �G��t<��t���_  �G0����H� �Y   H��0��G0����H� �   H��0��1 �G0   H� �   H��0���O8�  ��  �G0   �G    �   H� �s,1�A�   ��$  ��uJ�{��   �C�$�@�B H�C H��H�@h    �$�  H�{ �Y   H��0�<�C0    �C8  �   ����   �C��t}��tx�C0   H�{ �   H��0[�+����W(�w,1�A�   H� A�   ��#  ��u<�K��w4�   H��Ju�!t$�C4�C0    �C8�H�C H��H�@h    [�u�  [��AWI�   ����AVI��AUA��ATA���US1�QD��L���D�  A�ą��0  Ic�H��H-A�% H�}h u�1Ҿ   �@   ��d H��H����  H�]hH�C)�@ H�k D�k�C4�   �C,   A����   D���$ŀ�B H���]�  H�{ L�{,�Y   -   �C(H��0�   H���7�  H�{ �C0����-   �C(H��0��E�C0����H�}0�C(�   �[�C0   H�����  �C,   -   �C(;Et=H�{ �X   H��0�)�C0   H���ţ  -   �C(;EtH�{ �   H��0�2/ �   ����Z��[]A\A]A^A_�H���   H����   f�W�J�f��&��   �   APH��H�      H��u�   H��%H��uB�   H��#H��u�Y�xP uS�x\ uMHǀ�   ��B �0�xX u:�xd u4Hǀ�   �B ��xT u!�x` uHǀ�   �B �"   1��m. 1�Z�Y�����1��f�WH���   �J�f����   �   H��H��@�ƄuQ��  u'��AtpH����  �xP ua�x\ u[Hǀ�   E�B �BH����  �xT u?�x` u9Hǀ�   k�B � H����  �xX u�xd uHǀ�   ��B �"   1��- ATI��USH�O Hk�H*�% H�iH�]hH��tpf��f��}f���f��uuX�{0�u�C0   �(  H���  H�CH=)�@ t%H=�-A u�C,������   H�5��$ ���B ��J���C0������   H�}0f��t~��u�X   f��v�   �- 1Ҿ   �@   �a H��H��諲  H�]hH�   �   H�C0fA�D$H�C)�@ H�k �C,   f��"f��}<f��t-f��~P��f��v�Ef��ut1f��vu9�C   fA�D$  �!�C    ��C   fA�D$  ��C   �C,   H�����  -   �C([]A\��UH��1Ҿ   S�@   P��` H��H����  H�]hf�E  H�C)�@ H�k �C    H�C,   �C8  Z[]�UH��1Ҿ   S�@   P�` H��H��菱  �  H�]hH��H��f�E  H�k H�C)�@ �C   H�C,��  -   �C(H��   )  H�C4Z[]ø   ���   ��   ���   �u|H���   �zX to�wD��# DB@��+�% ����1�)�A9�|K�W��+�% A��A��D1�D)�A9�|.PH�Gp    �glH�=��% �A  H���% �zl��Z�����Ë��$ �F9WXu	9G��   AUE1�ATU��SH��Q�GH���% �WXH�GD9kp~jH�CxN�$�A�D$tUL���bO  �=�%  ~DI�D$H��% Hk�H�|H9�uI�D$ Hk�H�|A�D$@t�   ��u	����^���I���X[]A\A]��H�FX��$ 1�H�=�% H�8�5���USQH���   H��u1��?H���u+w�}+{�eJ  H���   �R@����+ 9�|�H���   H�����  ������Z[]�UH��SQH���   �ؚ  ��u1���   ���   �@t�࿉��   �   ��   ���    u�H���   �u�}+p+x��I  H���   ��  @��y( t��  �����   ������u
���  ~4눃�u���   �w������Ӂ��   1��H���t��u���Ӂ��   )���   ~����   D����   ����9����������   ��   E���Z[]�ATUS���   ��u1���   H����v���B 1��j���H���   H�ߋp<Hc��   ���Ze ��S�4� [e s�@  ���ŋ��   ��   ��s5�=��%  t,�S ;b�% ��  ��}��       �K �   ���   �k�=�%  �\���ǃ�      A�   ��% �B���% ��t;H�1�H��H�4ŠIf �@�  ��AE��щ½   �����������   r�C`�C ��[]A\�SH���������t����������   �   [�AWAVAUATUSH��H��H���    u��B 1��3������   H���   D�$�@[e �i�D$�A+CA��+k=  
 =  ��}fA�   �E1���  ��}A�   �A�   ��  
 ~_A�   ��1�����E�����H��� [e ���   D9�t3H���$�����t'�r  ��  ���U  A�   ��  
 A�   EN������=�   #��D������1�)�D��1�)�9�	D��E��A��E9���   E9���   A��tD���   H����������   A��u	�|$u�2D���   H���}�����t���   �D$H�߉��   �b�������   �2����   �tA1�����   H���:�������   �Ń�t'A9�t��܉��   H��������ui�̓��tA9�t���A��uǃ�      �ID���   H���������t��4A�   A�������3���E9��$����%���A�   A�   ����H��[]A\A]A^A_�AWAVA�����AUA��ATUSH��H�����   �h�1����l$Lc��   D�`B�<��9f  ��   D;|$��   ����   Ii�H  ��<f  ��   H���;f H����  ��tmH���;f E��tMi�H  I���;f H���   �   �`�P�H�s�{��  D��+S8����w�H���;f �p�x+s+{��D  =  @ ~��A�ċ��   �������   D���%���1�H��[]A\A]A^A_Ã��   �H��% H=`if t,H�x"A uH9�t���   9��   u	���    %H�@��H��h�   H�|$f�D$$��=���H��h��SH�GXH��Ǉ�       H� H�pH��u1�H���^�����u�   ���   t�H���   ���    uH���   �p��u�T茔  ��t����$|,��&~��("�����   ����r'��r����   ����r$���   H�߃����u1��# H���   H��[�p��N  [�S���   H����t�ȉ��   ���   H���   ��t"H��t	���    ǃ�       ��ȉ��   ���   ��&�C8��%   ���)υ�~-    �	��    EƉC8H��t	���   u!�   H���.������X  H���   �p�n���   ��t+$�=�r% ���   �-  �=�_%  �   H��[����H���   �x( t5H���������t)H���   �p��tH����! H���   �p(H��[��M  H���   �x, tH�=fr% �=�_%  u	���    u-H���������t!H���   H�ߋp,�M  ���   �   �   �=�h%  u
���   y1�;���    u�H���   H��舒  ��uھ   H��������t��>H��������uH������H���   �xP t�]�����H���   H��[�pP�! [�H���   H��tIUSH��R�w���   ߋH�P����  �C8H���   ���   t�����������)���k8X[]��H���    ttAUATUSH��P����D�k8�   H��D���>  H�߾   A���y  ����������)������   ��AY�D�H��[����D��]A\A]��D�R�   �n>  �H���    ��   AW�   A�   AVAUATA�   USH��R�  H�������D�k8�   H��D���y=  A������������)��
�����D��H�ߙD�A������D�R�   ��=  A��u�X[]A\A]A^A_��H���    ttAU�   ATUSH��P� H���m���D�k8H�ߺ   D����<  A������������)������   ��AY�D�H��[����D��]A\A]��D�R�   �W=  �SH�������I�����'~4H���   H��uH���   H��[�p��J  ���    ~�H����  ��t�[�SH�������� �����	~4H���   H��uH���   H��[�p�J  ���    ~�H��蹏  ��t�[�H���    tSH���o���H���   H��[�$   �V  �H���    t\SH���F���H���/�����t2H�߾7   �9 �k����   H���   H�ޙ���RH��[��"  H���   H�ߺ   [�RV  �H���    t>SH�������H���������t'�����
   H���   H�ޙ����   H��[�|"  [��H���    tOSH������H��������t%������   H���   H�ޙ����k�
H��[�5"  H���   H�ߺ    [�U  �H���    tSH���<���H���   H��[�!   �U  �H���    tTSH��������t2H�߾7   � �@����   H���   H�ޙ����k�
H��[�!  H���   H�ߺ   [�'U  �H���    tGSH�������C    �   H��H���   ��T  �k    �PpP�PtPH���   H���   [���aY% �R  ATUSH���W �w��
S  �S �   �s�{+st+{p�rF  �@x   H���n������   �   ��)��ȅ�N��   H���   H����   ���    ��   �U�M�s�{���  �S89�t1�Ƌ4�$ )ց�   �v��)�)��I��ʉ�)с�   �GЉS8D�c8H���$ A��B�4�H���   �x<�����B�4���B �CpH���   �x<������u�}+s+{�Ct��;  H���   �sx��y<�U �   ��  ( +S ��OȉЙ����    �� ���9�NщSx[]A\��H���    tSH������H�߾8   [�  �H���    t]SH��H�������H���������t>����H�߾5   �D$�� �D$�
   H��H���   H�������k�H��[�b  H��[��AWAVAUATUH��SQHc��   ���4  H���   �� [e H�=+r% �@<��W���Ze G�!r% �r% +�% +�% D��  ��D��  @ D��  ����  @ A��A��A����E9���   E��A9���   ���@ D��D����@  ����   H��q% H���   H��H���   ����H���   H��
  �E  H�=hq% �   � H�=Wq% H���   �sX�nE  �STH�>q% ���   �S�`l���   Hǀ�       Z[]A\A]A^A_�A���K���A���7���XH��[]A\A]A^A_�/����6   �( AUATUSQH���   H��tH��H���   �,Q  H��H��� �  ��taD�e8H���>  H��$ D�m�   A��B�4�����B�4���B �   D�D�m�C����H��AŋE D�k�C Z[]A\A]�a>  X[]A\A]�S�\   H��� H��[�O���S�[   H���i H��[�8���H���    tGSH���A���H���   �   �x�P ���`B  H���   H��H���   H���   H���   [������H���    ��   AUATUSH��V�����H���   H����  ����   �R   H���� �   H��H��H���   �z  H���   �  �L���   �H���   �~H�AxM��tf�k8D�i�   H���$ ����Hc�4������4���B �   A)�H���   E�l$D�h����H��L��F   A)�E�l$Y[]A\A]�!6  X[]A\A]��SH������H�߾c   [�
 USH��P������C8   H���   �O  H�ߺ	   H��H���,O  H��H�ߺ	   �O  H�ŋ@8��   H�Ų$ �]8����Hcۋ4�H���   �x<�����4���B �EpH���   �x<�ѿ���EtZ[]�USH��P�b����k8   H���   �N  H�ߺ	   H��H���N  H��H�ߺ	   �N  H�ŋ@8��   �H�4�$ �]8����Hcۋ4�H���   �x<�Y����4���B �EpH���   �x<�@����EtZ[]�AUATI��USP�����I��$�   ��M  L��	   H��I���N  H�ŋ@8��   �H���$ �]8����Hcۋ4�H���   �x<�ھ���4���B �EpH���   �x<�����L��L��	   �Et�M  H�ŋ@8��   H�Y�$ �]8����Hcۋ4�H���   �x<�~����4���B �EpH���   �x<�e����EtZ[]A\A]�ATUSL���   M����   H���   H�����      �p�� H��������k8�   H�Ѱ$ ���4������4���B �   �Cp�����A�t$A�|$+s+{�Ct��4  �   =�� ~
�   �����A�D$l��AD$ +C ����Cx[]A\�H�S�% 1�H=`if tH�x"A u���   u��H�@�݃���   AV�M�# �   AUATI��U��SH���   ��D�oB@�@�����   H���$ �ߋ4��1����4���B ��E�t$A�����A�L$ D��A�4��   �   ��=  �P�pH��H����+  ��uL��L��H�߹'  []A\A]A^�B  I��$�   H��H���   []A\A]A^�V����H���    tSH���?����s8H��[������S�G8H�����   ���   @������C8H�ߍ�   ������C8H��[��   �����SH���   H���p8��=��;}��tB�'��?"�����   ����r>�������   ����r;���   H�߃����u1�[� [þ   � H���   �p$��t� Ã��   ��H���   ��   �b1  �5��# ��b% ��u����  ���   ����   ���$�=��# ���   w���^  ��ut�=�Z% �L  �e��Z% ��t��uC��A�����"��t��t#�+��A�����
��A��������D!����u�������������   1��<��9f  tHi�H  ��<f  
H��H��u��H�~�% H=`if t0H�x"A u H9�t���   9��   u���    ��   H�@��H��h��u#��uh���   ��t-��uXf�D$$��   �&��Y% ��t��u:��t��u0f�D$$��   H�|$�  ��   H�|$f�D$$��D�����,���H��h��S�T   H��� H��[����S�U   H��� H��[����S�O   H��� H��[�~���H�?�   �t H�?�   �g UH���   SH��PH�?�Q ZH��H��[]�R  ��g%     H�1�% 1�1���%     H=`if t(H�x"A u���   uHc���H��`Hf �H�@�Є�t��g% �`   1��� �a   1��� AUI��ATU�   SR�G��  <�A�E��?9�|nA�ED��  ��������!   D��������   �9  I�������  L����	A�D$x�M;  ����A��$�   ��)��ɉ�NŁ�   A��$�   �X�b   [1�]A\A]�, ATUH��SD�g�S������L����m)��B������!   ��D������   ���9  H������H�߾  ��	�Cx�:  �������   �   ��)��ȅ�N��   []A\������H% ���=,_% �6% ��thUSH��PHc% H��H�,�`Hf ���H���=f% �% �   �F  1�H���   H���E+CH���   ��yt��~�^   ���   Z[]�! ����   ��   UH��SRH���   �(F  �   �P �pH�Ëx�8  �#   H���� �����   ��1~j�   ��Y~`�   ��w~V�   =�   ~J�   =�   ~>�   =�   ~2�   =�   ~&�   =�   ~�   =�   ~1�=�   ���L	�s�{�S �7  �   H��H��������tH���   H�ߋp�9  �S�sH���N"  XH��[]�p8  �S�_   H���
 H��[������=�{# �9   u1����   �@�ƃ�9�� ATU��SH��E��t
A��tr��   A���t
A��t$��   D�'D��)�9�|����!,  ����   �9D�'D�9�~���H���,  ����   D�#�}�7����+  ����   ��t@D�#�1A���tA��t7�pD�gD��)�9�|3�G���+  ��uU��tD�c��H���+  �   �=D�gD�9�~&�S��H���+  ��uD�c��H���m+  �   ��w���\+  1�[]A\�UE1�SH��Q�O�W4�w8D�K(H� ����������% uH�C �   H�x0� ��uOH�C �S(H�@h    ��u�{���u�{u�S,f�P�S0f�PH���=�  H�{ �   Z[]H��0�E X[]�AW�    AVAUA�   ATA��USH����	AD�H�<$1����D$H�<$����  �Å��  Lc�M��I��L�z% I�xh M��u�1Ҿ   �@   �? I��H��芐  M�uhI�F��@ E�fA�F    A����  D���$�8�B A�F(����L��M�n A�F8   �!~  �  A�F(����L��M�n A�F8   ��}  ��   A�F(����L��M�n A�F8   ��}  A�F4A;E �(     �   A�F   A�F(   L��M�n A�F8   �s~  A�U9�O�A�F4�D$A)F4��  A�F(   M�n A�F8   �A�F(   M�n A�F8   A�u L���}  �<A�E A�F(   M�n A�F8      �A�E A�F(   M�n A�F8      A�F4�c  A�E A�F(   M�n    A�F8   A�F4H�$H�@8�Pf�@fA�UfA�E�$  A�F(   A����1�M�n A�F8   A9mp~`����7|  ��tO1҉����{  H�@
f��xH���% ��A9�DO��   ����{  H�@
f��xH�|�% ��A9�DO����I�F D8E�~4�   A�F(����L��1�M�n A�F8   ��{  A�F4A�EfA�F0A9mp~a����{  ��tP1҉���'{  �   H�@H+5x% H��L9�t1҉���1{  I��A�F4A9E uA�EfA�F0A�EA�F,���뙽   �����H����[]A\A]A^A_�AWE1�AVE1�AUA��ATE1�U���SH��(H�<$H�<$���|  �Ņ��U  Hc�H��H�w% H�{h u�1Ҿ   �@   �K< I��H���H�  L�shI�F��@ A�F(   I�^ E��tA���   DD��   DD��A� @  A�   D�D�[E�~8E�E�N4A�   �spL�w% 1�9��M���H�CxH���A��   H�A8L)�H��9���   H�I@fD;YuE�H�yh uu1Ҿ   �@   H�L$D�L$L�T$D�\$�t; H��H���q�  H�L$L�T$D�L$D�\$H��H�YhL)�H�C��@ �C(   H��H�K D�{8D�K4H���=���H���A���H��(D��[]A\A]A^A_Ã��%  ATA��U��SH����v���B 1��������H�<����   ���   9�u1���   ��p[e E��tA���
A�   �A���{V% ����u��9�L����   �   ����   ��t?��t��tV��tq�   �{| �   u���    tǃ�      �jǃ�      �^�{|�   wS���    tJǃ�      �>�{|�   w3���    t*ǃ�      ��{| �   u���    t
ǃ�      []A\�1��AUATU��SI��H��Q�=}L%  ��   ��M% ��t{��uwH��D���   E��tE1��   Hk����   ǂ�      �   ���_d ��u�   H���[���Hc�J% D���   Hi�H  H�;f H9�u��!   1��| �WHk����_d 1���t��t�   ��   H������H��1҃��    uǁ�      �   D���   E1�	�A��ZD��[]A\A]ËW,1���c�d   H���dO։W,���   �   �k�d1�9W0}�w4�   �W0É�H���xP uǇ�      �@P   Å�u	�G8  �e��uH��G@4  ���      �J��u	�GLh  �<��u	�GD4  �.��u�d   �P����G<   �Hc�1�H���z8 u�B8   �   ËG +F 9Fl�B  =  ���7  ���    �*  ATI��US�G<H���   ��7��&��  �$�x�B �{0c��  Hǃ�   ��B �  @H��H�C0�  �{0�   ��  Hǃ�   ͬB �  @H��H�C0�e  �C,��   ��=�   O�H��C,���   Hǃ�   �B �7  �C0��   ��=�   O{4 �C0u�C4   Hǃ�    �B �  �C,��   ��d=�   O�H��C,���   Hǃ�   �B ��  �=�p# �  H��C,�   �   H��ǀ�   �   �����Hǃ�   '�B ��  �{P uHǃ�   3�B 1�H��������=/I%  ��  �k  �{T uHǃ�   M�B �   �΃{X uHǃ�   i�B �   붃{\ uHǃ�   ��B �   랃{` uHǃ�   ��B �   놃{d uHǃ�   ��B �   �k����
   H���������&  Hǃ�   ׭B ��  �   H����������  �{,Hǃ�   �B �  Hǃ�   �B �  �C8  Hǃ�   ,�B �   �d   H�߽]   �����{| �C<   Hǃ�   =�B �P  ǃ�       �A  H��C@4  ���      Hǃ�   F�B �D�CD4  Hǃ�   [�B �0�{H �H  �CH   Hǃ�   t�B ��CLh  Hǃ�   ��B �]   ��  �   ���   t1�1�H����������  Hǃ�   ��B �  1��   H����������  Hǃ�   ��B �t  �   �   H���W�������  Hǃ�   ήB �J  �   �   H���-������{  Hǃ�   �B �   �   �   H���������Q  Hǃ�   ��B ��  �   �   H����������'  Hǃ�   �B ��  �   �   H����������  Hǃ�   7�B �  �   �   H����������  Hǃ�   S�B �x  �{h u1�Ѥ�   H��H��u��Ch   1��   H�����:�����u�Hǃ�   v�B �0  1Ҿ   H���G������d  Hǃ�   ��B ��   ���   �   H�������������3  Hǃ�   ��B ��   1Ҿ   H����������  Hǃ�   ίB �   1Ҿ   H�����������   Hǃ�   �B �z1Ҿ   H����������   Hǃ�   �B �V���   �   H�������v�������   Hǃ�    �B �(���   �   H�������H�����tiHǃ�   5�B �!   ��P�B 1������    A��$�   �t���   L���{(  HctC% ���   Hi�H  H�;f H9�u[��1�]A\���  []A\��S���   H����������   ���   t%�������   ���   �{l��  H�����   H���   tCH���   H��t7��s���   H����   I�������H��H���;f H��I���D�l��=�C%  u��s��H% H��tnH��u H�������H��H���;f H��H���D�l���H�ǁ�  ���   �@   �f=  HcRB% Hi�H  H�;f H9��   u�=՟$  t�*"��H���   �P��9��   }�p4��u�p0H���'  ��������   �   ��)ǅ���N=j# 	���   tH���   ��tw�����
t��u-�?   ��M   ��I   �s�{�   ��t%  ���      [Ë��   ���  AWAVAUATUSH��H�����    ��  ��I��I�Չ�sH�Gp    �Gx    L���   M����  �=sK%  u��M����   ����   M��tI���   H��t
�x|��   �K�SL�D$A�pA�x若  H���   A��i� � ��yHA�ǃ�'/9��   }'L�D$�C A+@ =  @ ~�����tA��   �A��H�O�$ A��D��B�4�聣��CpB�4���B D���n���CtM����   H�CXH� f�xu���   9��h����  A��$�   ��  A�|$8 ��  A�D$4��t0�ȹ   t�   ����A�T$09�A�D$4    ��)�)�A�T$0A�D$,�    M��$�   )�Hºd   A�D$,A��$�   ��dO�A��$�   Hc�?% Hi�H  H�;f I9�u��d�
   �(   NՍT(�Y������   )艃�   ��H��H��L��[]A\A]A^A_�����6���H���   ;B } ���   ��r��@�rH�߉��   �$  ���    ǃ�       t	���   unM��tiL9�tdA���   tZH���   L���   ǃ�   d   HcBHk�(H �d H9��   u+�r��t$H��H��[]A\A]A^A_�<$  M����������H��[]A\A]A^A_���O u%H�G�W$�H9�u�W(f�P�G0�f�P�G,�G ËG(���t��t!�H�W�J�A�f�B�;G +f�J�G(   �H�W�J�Af�B�;G$|f�J�G(������O u4SH�������H�s�����N�C(��)�9�|�C$)�f�F�C    [���O u7H�G�W$SH���H9�u�W(f�P����#C0�f�P����#C,���C [��UH��1Ҿ   SPf�G  �0   ��+ H��H����|  �uH�kH��H�C��@ �s$�l  �C    ���C(Z[]�UH��1Ҿ   SPf�G  �8   �+ H��H���|  �uH�kH��H�C��@ �s$��k  �C(�  H��H�C,�����#C,���C Z[]�AUA���   ATA��1�UH���8   SQ�.+ H��H���+|  �uH�kH��D�k,�C0   H�C0�@ �s(�Uk  �C$;C(u�C$    f�E  E��u�X��������C ��C    X[]A\A]�UH��S���R��H����j  �Å�x#Hc�H��H=�e% H�h u�1Ҿ#   �<�����X[]�AVI��AUE1�ATUSH��e% D9-�e% ~GA�Ff9Cu4�kE1�D9cp~#H�CxH��J�<���h  H��t	�@9�O�I����f�kA��H���[]A\A]A^�AVI��AUE1�ATU��SH�:e% D9-Ce% ~GA�Ff9Cu4��u,E1�D9cp~#H�CxH��J�<��mh  H��t	�@9�L�I����f�kA��H���[]A\A]A^�UH��1Ҿ   S�0   P�) H��H���z  H�k�uH����i  �C �EH�C[�@ �C$�C(����f�E  Z[]�S�   H�����   ����  �G+�M% A��H�5@N% A��D1��NhOhD)�9��x  �G+WM% A��A��D1�D)�9��U  H9��L  ���   ��shH�|$�K����   H�|$H�5�M% ���H���   �JH���HL����H�=�M% H���   H�Gp    ���   �����Gx    �p�  �   ����   �O D�Gl�   �F A�D9���   Fl9���   H���   H��t4���   ���   9�t��u��t
��u��u�   H9�ts1ۅ�um��u
1ۀ����^H�|$�d����   H�|$H�5�L% ���H���   �JH���   �HL�����1��"1����À�t�M% t������   H����[�UH��SQ� u���B 1�菋��H�]�CuIH��L% H�ڋp�x�.  ��uh�E ��L% 9�}b��L% H��L% ��L% H�fK% H�L% �?H���/  H�6L% �Hl;�L% ��P ��L% )�9����L% )�=   ��   �1�Z[]�AUATI��USQ�oH�_����   �Cu1��5  H����  �dL% 9jL% }�A�4$�=�K% �'�����H�C@H��t
H�S8� 9t!�=>L% ��+=�K% ����9b% }�b% H�C@H��tH�S8�@9Bt!�=�K% ��+=�K% �ۚ��9�a% ~��a% 1��a% 9�a% @���   H9;K% u�   �}���   t��7�=K% �~����{l{ ��+=VK% A���z���9ta% A��{ D��+=7K% �^����La% 9�|�9Na% MGa% D9�   AO�H�(K% Й����I% Z��[]A\A]�AWAVAUATUH��SQD�gH�_E���r  f�{ tH�=~J% H���i  �Cu~�5bJ% �m �   �љ���=�V% D�%�V% )ŉ�詙���=�V% ��D�-�V% A��蒙���5"J% ��A��肙���=6I% ���u���H�K8QJ% ���A
;=�( ��   ��   H����  �u �=�I% �>���A��H�C@H��u"�=^J% D��+=	J% �0���9�H% �@����FH�S8� 9uH�C@H�S8�@9Bu,A�   �  �=J% D��+=�I% ����9�H% }�������=�I% D��+=�I% �Ș��9jH% ������9Q|H�K@H��t�I
9�tC�t= C�<4��%  E1��  H9I% �y������   �l����7�=�H% �U����{l{ ��+=-I% A���Q���9�G% �=����{ D��+=I% �4���9�G% � ����5�H% D�m �  
 �����=*U% D�5U% A)�D�������=U% D��D�=U% A��җ���5bH% D��A�������=uG% ��贗���H% ��H�E���   tD��D����$  ���H% D��D���c%  �yH% �������H�5
H% H��H�������ZD��[]A\A]A^A_ø   ���   tm�G+G% �H�5�G% 1�)ЋNhOh�¸   9�~G�G+�F% �1�)�9�~/H9�t*H���    u1��=B>% uPH��'  �W����   Zø   �ËG,9�G% ��  �G09|G% ��  �G(9eG% ��  �G$9ZG% �u  SH��H���pJf �9  ���U  1�H�{@ �M  H��F% ���   u�S���1  H���    u	���  H���  �]G% ;�F% }��F% H�8G% �NG% ;�F% ~��F% �S% ;�F% }��F% f�{ ��   Hc�F% H��H�ՠIf ���{F% ����   �=�$  u7�   �ϱB �ω����~H�@% H���e H�|�������
���$ ���H+\% �%F% H��i�z�E��$ ��t#��	|$��	Hc҉�pJf �(��u�3F% ��E% �H�=^�$ �رB 1��R	���   [ø   �SH�Wf�z u)H���  �=BF%  �   AH�=�E% �Q   ��  �,H��E% H���p�x�  1�H�sH�=�E% ������l  1�[����   ��   ���   �����trUSQH�5CD% �G�_+F+^�1�)Љ���1�)�9�M�+_h�    ��H�9tE% ~*H���,\  ��t�`E% H�=E% H��H�5�C% )�����Z�   []ø   �AW��A��AVI��AUATUSH�����   ��C% �T$��D% �Gh�5�C% �H�=oD% D����D% �ʉ�)�)���D% �0�t$��D% �}D% ��  �rD% �-pD% H��D%     H� D�%SD% D�-HD% ��@�)D%     ��\$ �D% ��Y% �ED% )�)ŋ�Y% �1D% ��    ��    ��A)�A)���A��    A��    A��A��9�.E��E9�"�hA D�Ɖ�D�D$�  ��tCD�D$A��������L����  ��C% E�~L��A�F`�vC% A�Fd�D$A�F�E  �   H��[]A\A]A^A_�AV��AUATUS���   �5gB% �yC% �OhH�=C% �Ǎ4)ωBB% �54C% ��)Ή=2C% �ǉ5&C% �4�5%C% ��軙  H�gC%     H� ��@��B%     ��[$ �C% �C% ��B% ��B% ��   ��X% ��B% �-�B% ��X% )�D�%�B% )ŋ�B% ��    A)ԁ�    ��)�A��    ��-    A����A��9�|(E��E9�|���@ D�����X  ��u1��uA�������ԋ X% �JB% D�%GB% D�-8B% )Ë-,B% A)ċ�W% ��A��A)�)�A����A9�|$E��D9�|��A D�����p  ��t�A�������׸   []A\A]A^�AWAVA��AUATU��SH��Q��A%     �J�����u1��,  ���   ��sPH���  D�cD�k�k��A% D�sH��I���.�袋.�C`�QA% �Cd�)  ���    �  ��   �   �.A% �dA% �{l��)�9�|��gA%    ��r�s )�9��i�����)��   �Y�����D�c���+!A% =   �R����:���H��s�{H�,ŠIf H���b  H��D��D��A���Q  A9�u��@% �B���@% ��u��   �%f�} t�H��H+=\V% H�ډ�H��I����[  ��Z[]A\A]A^A_�ATUS�WH���wD�g �o`������u@% �3@% �S`�CdA9�u�S ��Kl�s �9�}��)ω{ )�;Cl[��]A\���USH��Q��������   ���    !�  H����  ���   �H�Ch    �   ���   ��s
H���  �|�tx�=�>%  ��?%    te��^% u\H�߹
   1�1��U����Cl�   �s�{����&   C ���  H��蠯����虯��)����]p茯����腯��)����]tZ�   []ËG4��u�3>%     ���u��?%     �H��>% ATUSH���p�xH���  �K�S1�A��1���  A�̉�u��   ���=% �D?% 1�1��ŏ  )��=   �v��   ��5�=% �=?% �����  H���$ �ǋ4�����A��H���$ D��4��ύ���4���B D���>% 躍��[]�h=% A\�AWAVA� �  AUA�   ATUSH��H��H�=>% A��u8�s�StH��S�R�������  �sp�SH��sH��[]A\A]A^A_�+���D�c�kh�SpE��A�A)��	D��E��A�C�KtA��A)�Ņ���D��A���D�A���@ ��A�   D��D�T$��=%   �c  D�T$�Kt��SpA���@ A�   D���D��=  �Kt�SpD��A���@ A�   D��D�D��  �5}=% ��  �	�����   �5e=% ��&D��+5X=% �   ��   O��5D=% ��8�   �{p�Q����{t�5*=% ���A����sCH�߉��������u������{p�����5�<% �{t�-=% �
���H�=�<% ��;% �j����5=% ��;% H�߉sps�StS�������E���H��[]A\A]A^A_�U��S��Q���  A�؉�A�H�@ ���x�pH�5<% H�N~$ B���-<% ��R%  �  ��R%  `����B����B D�@lH�]<%     A��D@ ��A��   ��D�"<% A�   �	  H�=/<%  ��:% u1�Z[]���D�<% ��I��A��H�5�}$ ��H�=�;% �F��A�q�};% ��:% D��B����B A�   A�D�0A�AlD��D����AA A���@    ��;% �	  H�A��A A�   �B8�zH�S;% �r��HcЉ�����B H�*}$ ����������  AV�ы�P% AU��D��P% ATUS�_H�=�9% D�$)�H�5;% A)�)ËG�-;% A����D�,)ȉ�E)�D)�A����D9� A��E9�D��� A ��A���  ������[]A\A]A^���:%     �5�9% ATUH��S�_(9],|"D�e$D9e |D��T
A ��A���E  ������[�s:% ]A\É�E1�1�Hk�Hc׋�@�B ��t[D�H��9�~LHk�H��H�B H��@�B H��t:D)��z tA�   �A��H�H�f�4��f�t�A�   �A��H��4��A���Á�   I��6Dk�D���u���A�rA�y�h���I�rA�y�[�������1�)ǉ���1�)ƍ79�}��)����)�ËB�JL���u����A;8U���E�H��uA9�|��Å������ATD)���U��SA+8H�Ӊ����m����s��A���_���[]A9�A\������ATUS�F4��tP��tI��H����ts����   1�1��   H��~ ��W�@x1�9�@��9����-1�9�@��9����H��~ �O�W� x1�9�@��9������C1�9�@��9�����H��3������s�{����H��3������s�{��L�������9�t���[]A\ËBD�B��uD����9:|tE���D�JE��uD9���Å������D1���+
D)�1�AT1�U��Sy
��D1����/��D��H�Ӊ��������s����A��������A9�����[]A\��H���@�F�G��F�G�F�AUI��ATUSH��AP�w�{������{A�u����豆��)�t8�s�;A+} ��蜆���sA�}+{A����臆��Y��[A�<]A\A]釆��Z1�[]A\A]�USH��H����C%    =    w�|C%    =    v)H���Vf �p�8������Vf ��H�C�p�8�����6H���56C% �=,C% �D����5-C% �=#C% H��5C% =C% ���"���9�tlH��H�������H���Vf �������xP�=�6%  t=��  	1�H�{@ t<H�5�6% H���H�� Kf �F   H��H�^���   ~�f���H��6% �   H����[]�AWAVAUI��ATUSH��(�oh�G�_A���A��A)�D$�A)�[B% 3YB% ~D��A�܉ú�Vf D��D�������|$��Vf ��A���x���A9�ta�D)�H�t$��Vf D�t$D�d$�l$�\$�������x7H�5�5% H���H�� Kf �F    H��L�n���   ~����H��5% H��(�   []A\A]A^A_�f� �u��5%     �H�W8H�O@�A�	9BNB��x5% 9�~�z5% �XA% ��l5% �JA% +`5% �f5% Ë��   ��u+H�G(H��tH�O0H�H0H�O0H��tH�A(�H�OXH�	H�A`��ueH�wHH��tH�GPH�FPH�GPH��tH�pHËG+RJ% ����x6�G+>J% �����[J% 9�~��x9aJ% ~���H�[J% H�H�4��SH���w��֊  ���   H�CX��u H�H�C0    H�A`H�C(H��tH�X0H�Y`��us�C+�I% ����xS�C+�I% ������I% 9�~;��x79�I% ~/��H�CP    �H��I% H�H��H�H�CHH��tH�XPH��H�CP    H�CH    [Å�xs��xo�rI% 9�~e95|I% ~]��UH��SQH�:I% �H�H�BH�H�H% H�;f���u�   �%Hk�XH=�H% ��K$ 9GHuH���ӉGH�Յ�u�Z[]ø   Å�xM��xI��H% 9�~?95�H% ~7��UH��SQH��H% �H�H��H��u�   �H���Յ�tH�[H��Z[]ø   �AUI��ATE1�U��SQH�3% H�� Kf H����tAH�53% � Kf ����H9�v�9�}I�ĉ�H����9�L����A�Յ�tA�$���뻸   Z[]A\A]�AWD��AV��AUATUSH��8��2% ��D�D$D��G% L�L$ D)���J$ H�|2%  Kf ��� u��   ��G% A��A)�A���� u��   A�։�D)�)�A)�)�=/>% D)ǉ5*>% ��)����������T$��A��D�5>% A���	>% A���t$�L$(9�}.��A�   ��A)�D������D1�)�蹀���D$   �D$�>~&D��D��������D1�)�葀���D$�����D$��D$    A�   �D$   �t$D�����L���D�| D;l$(}'�Ž   D��A�   )ŉ���1É�)��/������-~��D����A�����1É�)��������E1��   �   ��޽@   ����AċD$���D$,�|$, u	�D$t.��|$�OA D���������u��s�|$�YA D���G�����t^�T$9T$uD9l$(t0D����D9�u�L$D|$L$�D����;D$uA�E���u�H�|$ H��8�   []A\A]A^A_�<���H��81�[]A\A]A^A_�AVA����   AUA���   ATA��U��1�S�m
 �8   H��1�H���Ik�\D���   D�sD�kH�jd �=&% �P@H���   �Sh�PD�Sl�PT���   �P���   t	�@���   胟���   Ik�\H�ߙ��Hc��jd Hk�(��(�d ���   ���   H�� �d �� �d H���   �C<�B�C@�����H�CXH� ��@�S`�Cd��   �u�S ������uH���   +BD�C ��k H�C"A H���zZ  H��[]A\A]A^�S���   H��%  ��ub���   �����8tTHc8B% H���   Hk�
H������;�:% H�� Yf ���   �B% f��(Yf �/M% �� Wf u������:% H���V���H�����  H��[��Y  USH��Q��uHǃ�       H���U���1��U��Hk�(H�� �d ��(�d �� �d H���   �S<�PH�@���   �S@H��tH����Hk�(���    ��8�d t��   Z[]�S���   H��H�Gp    Hk�\�Gx    ��kd �^���諝�����   �   ��)��ɉ�N��   �������   H���   �p8��t	H��[�6�  [�USH��QH���   �G H��t�W`9�~�q )�)ֺ  ) )�q ���Q$���   Cx�C ��s\H���   H��tP��   uH�s�{+p+x�;���H���   �Sl�K ��V )�yk����   9��t�R9�~	��   �K �C`9C |�-A# ��v���   t�[x�Cx��y-H���   H��t=  ��}���"   H�߉B$�G�  �Cx    �C`�C ���   ��w	��s�[x%  =   u,ZH��[]�n������   u�Cx��u	�Cx  ���-   �Cx�Sl�K �Cd�9�~-�{x ~�Cx    )ЉC ���   ��s�[x%  =   t�X[]�H�p u1���   ���  %�����Gx    ���   H���   �p�[���AVAUATUS�GpL���   =   ~	�Gp   �=  ��}�Gp  ���Gt=   ~	�Gt   �=  ��}�Gt  ��D�gp�otH��A�   �s�KA��   ��   ~D��A���A��Ɖ����A����D�T E1�1�H���������u`H���    t
H���]����L���   t;H�+% H��t%H�@@H��t�@
;�g( uH��[]A\A]A^�����H��������H�Cp    D��	��M���M��tA���   ��   ���   �  ��   �S`9S ��   ���{ps'�� @  = �  w�Ct @  = �  vH�CXH� ;u���  =�  wU�Ct�  =�  wFM��t7fA�} u9I�} H���   H- �d H��i�����-�   ��w
��   ����H�Cp    �� �  ��x���{t� �  �Cp��x���Ct[]A\A]A^��ATUS���   H��D���   ��A����D�����������   H�CX�s�'   �{H� ��]����#   H���$�  D�����  �'   D���H� ��2����#   H�����  H���   1҉�   D��@T%   �������������-   H��H���   H���   ���   f���   f���   ��f��f�����A8���   t���    ǁ�      H��[]A\�����[]A\�SH�p H��u���   u
�C`9C t�'H������H�{�u��   �{x u���   ���u�.H�������H�{�u��`�ȉ��   uVH���   H��[�p��������   @t:�=�%  t1���   �����   =�  ~��F% u�������	H��[�9���[Ã=P% �$  AUATUSRHc,4% 9F;% �  �jF% +� Wf =  ��   Hk�
�� Yf D��"Yf L�� Yf ��A��D�����}  �(   D���H� ��^����Z   H���%�  A�U1�Hk�\��;��jd tH��H=�   u繉   Hc�1�D���Hk�\��4kd %   ����Hk�
�����������-   H�� Yf H��H���   f��(Yf f���   f��$Yf ��f��f�����A8�)3% �����3% X[]A\A]���Gf���>  ��ATUSHc؃<��9f  �"  Li�H  H��I���;f A�|$u���>���u�} 1ɺ   ������L���H��f�Ef��~��-   	��   f�E�-   L���   L���f��f�����A8Hi�H  H���;f �S,���   �C    ǃ�       Hǃ�       Hǀ�<f     Hǀ�<f     �C   ) H���;f �  �='%  t*�CP   �CT   �CX   �C\   �C`   �Cd   �E��;�% u�u�  []A\�Y��[]A\���wf��u*H��:% H=�_f ��  H�H�f�WH��:% 
f�P�f����  f��0��H�Hc�Hk�
�=�%  H�� `f f�Gf��`f �n  �A����=/%  �Wu	���S  �:% �   ��t��t������   ���,  U1�SH��RHk�\��;��jd t#H��H=�   u��K��h�B 1��$c����   �=�%  tHc�Hk�\��7kd ��   �= %  t����   Hc�Hk�\��6kd @��   Hc��;�s1�Hk�\������4kd %   �������� ���H��H����    H���   f�Cf���   ~��������   ���   ���   ��s�|% ��s�t% f�C�-   ��f��f�����E8�Ct	�� ���   X[]��U��SH���|$�t$�w������p����t$�|$�%   )���
�+�K����@x   H���G������   �   ��)��ɉ�N=�"%   @ ���   uH��H�߾_   []����H��[]�ATA��U��SH���|$�4$�����������4$�|$�&   )���
B�#�����@x   H�$躒��H�<$�   �[   �����   )��ȅ�N��   �E���v
���\   H��[]A\�#���H��[]A\�SH���c����   �spH�ߋ��   ��)��ɉ�NSt��s�s���   �Cx��S��C �S������u	H��[�;���[�H��H��u$H���$     � �e ���$     ��$     �AV��AUI��ATUH��S�G �w�    ������H��H���   �p��tH���o�  A�MA�UH���   �u�}�Nr  A��A���   t�z���A���r���A)�A��E�H�9c$ D�c8A��B�4�H���   �x<�`p��B�4���B �CpH���   �x<�Fp��A�uA�}+u+}�Ct�P���H���   H�ߙ�y<�   ��A�E +E ��Nʙ���Cx�~���H��[]A\A]A^�AV�   A��AUATI��US�o8�������H�=� %  A��uL��   �   L��������H�=� %  A��u*��   ��   L��������H�=� %  A��uA�\$8E1�A�D$ A�t$D��A�|$��    �>���H��H���   �p��tH�����  H�b$ �]8��L���   �4�H���   �x<�$o���4���B �EpH���   �x<�o��D��EtH���   �x<��n��H��Ex[]A\A]A^�]���1�H��@^f H��t9x@u�x4u�H8H�@�-A �H4H��H��u��1�H��@^f H��t#�H4��t�w9p@u�H8�@4   H�@    H��H��u��1�H�<�@^f  uH�H�<�@^f �H��H��u῕�B 1���]��AWA��AVA��AUATUH��SH����u	��A���A��1�A���D�|$D��H���9  A�Ņ���  Ic�H��H�4% H�yh I��u�1Ҿ   �H   �B�  H��H���?J  �ED�sDL�{I�_hH�C�-A �C<    �C@A���  D��M�g0�$��B H�EA�7�C  �  L��Hk�H�3% H�@�@fA�G��7  �C,    �C(�C4    fA�G  �;H�E�C  �  Hk�Hh3% H�@�@fA�G�D$A�C,    �C(�C4    �   �z�C    ��C    L���7  A��C,i   �C4   9ЉS(OC$�?�C    L����6  A�L��9�OC$�7  A��C,i   9�LC(�~������C4�   L���4�  H�߻   �����^���H����[]A\A]A^A_�S1�Hc�H9<�@^f uH�GH�@h    ��H  H��@^f     [�H��H��u˿��B 1�[�[��USH��V�G4����   ��t����   �  �W(�O<A�   E1��w H�诵���ŋCD�P���w�`;% uH�C�   H�x0�e�  ��u �{< ��   �C,H�{�C4   �C0�   ����   �C,�C4   �   �C0H�CH�x0��  �CD�ȃ�wlYH��[]������W$�w A���E1�H�1�������uD�C,H�{�   �C4   �C0H��0� �O0u#H��C$9�����C4H��0�   Z[]��  X[]�Hc�)���   �AULc�ATUH��SIk�QL��  ��uMk�JǄ-      �z��H�L Hk�(H �d �pH��  ��  �p��t�@ ����  ����   Hk�(H��0�d H��uH�D H��  ��   �Rt��L��H����H��   u�X[]A\A]�Pk�9% u�(%�  �4���B �j��k�9% u�ǉ�/% ��   ���  �4���B ��i���؉f/% Z�S���   
H��u	�G|���   ���   uH�;�
   �i�  ���   H��1�Hk����_d ǃ�   
   ǃ     � [�����W|Hk����_d �(   ��t
1Ƀ������   ���/  9���   �"  Q���    t!���    t�=o.#  tǇ�      ��   ���    t!���   ~�=E.# uǇ�      �   ���    t���    tǇ�      �   ���    t���    tǇ�      �y���    tǇ�      �d���    tǇ�      �O���    t���    tǇ�      �1���    t���   (~�=�-#  tǇ�      �
Ǉ�       Hk�1����_d �M���1�Z��SH��������t0H�;��   �����C|H��1�Hk����_d ����H�;[H���h���[ËG|1�Hk����_d �����ATI��USH��H�?H���   H=0�d tH=X�d u
��   �?����{|uI�<$��d uH�;�   �=�  ���   
u�{, u�C|H��1�[]A\Hk����_d �����Ct*���    t�C|�����t ǃ�      H��[]A\����ǃ�       �-�6% H��Y$ �{(�����  ��  �4��g���4���B �{(   A�D$��f��[]    A�D$A\��Gt���   
u�, t���   ����Ǉ�       ���������F   �F=�� ~+�u�F  � Ã, u	1�1��������   �G|����ËF-   =    ~�FËG|�F    1�Hk����_d �U���SH��H�?��   �����C|H�߾   [Hk����_d �)���ATUH��SH�������
   ����}< D�DtEk�
H�E D�D$D�`8躆����賆��H�} �  @ )���D�������D�D$H�} �މ��  @ ����H�=�%  t-H�} �S   �5�  H�] H��% �s�H�P�{�g  �C8H��[]A\�AUATUH��SQ�5���A��H�E D�h8�%���������H�} � @ )���D���_����
   H�} ��D�������D�D� @ �����H�=�%  uH�} �   Z[]A\A]鎻  H�} �   耻  H��% H�E �J�p�R�x�]f  H�M �ƋQ8)ց�   �v��333�0������M����333-�0��333FA8���   �   X[]A\A]�P�O|�   Hk����_d �\����!   H�?Z�E���P�O|�(   Hk����_d �6����#   H�?Z����U�   SH��P�G|Hk����_d �����G|Hk����_d �΄��H�߾   ���(�����H�;�"   Z[]�����UH��SR�_8�   �������H�=�%  �)% u<��   �   H�������H�=�%  ��(% u��   ��   H��������(% X[]�ATI��US��H���4����   A�l$8���D�BG����uD�D$�������
���D�D$)���݋�(% H����L��[�   ]A\�����SH��H�?�   虹  H�;��   �q����C|H�ߺ   Hk����_d ������C|�   Hk����_d �����H�;�����1�H�;���    @��[�.���U�   �   SH��RH�?�%�  H�;��   ������C|H�ߺ   Hk����_d �`����C|�   Hk����_d �T���H�;�k���H�;1��������u�X[]�AW�   AVA�   AUA�   ATUSH��RH�?覸  H�;��   �~����C|H�ߺ   Hk����_d ������C|�   Hk����_d �����H�;�����蒂��A��H�D�`8胂�����|���)��u�����D�A���g���H�;���D���A)̋�&% A��A��D���D���   �8���A��u�X[]A\A]A^A_�UH���   SH��QH�?�۷  �C|Hk����_d ����    ��   H�;��   �����C|H�ߺ   Hk����_d ������C|�   Hk�Hc��_d H���������Hk�(HU H��@�d H��H�������H�;�����1�H�;���    @��Z[]�1���X[]�Ǉ       �Ǉ      �Ǉ      �AUATUH��S1�R�E8H���   �   ��   �����H�D% H��tM�Pl�p�*   E1�xA�   ��P ������������E�dA��u�H���   H�=�% D��H���_����Ù�������?�z���X[]A\A]�H�?�	   �t�  HǇ      �G|HǇ(      ���   ����U1�SH��RHk�H��  H��t$��  ���t�ȉ�  u�Q��H������H��t�   �H��  H��4  X[]�H��H��$% �   �   @�|$H�|$����H��u$�=�$%  uH�53Y$ ��B �i�����$%    H���S��@��������[�S��@������������������@���w�����[�o���SH���?������{�����H�{[�SH��������{����H�{ H+=%%% H�������{(�����{,�����{0�|����{4�t����{8�l����{<�d����{@[�[���U1�SRH�=�#% ��������ۃ�9�t1����������X[]�H��H��#% �   �   H�|$�)���H��u$�=}#%  uH�5X$ �5�B �:����`#%    �D$H���S��������������	�[�ATUS����D���������}��������r�����	���[D	�	�]A\�U1�SRH�=�"% �'������ۃ�9�t	�?�������X[]�SH������H�H�����H�H�C����H�H�C[�H�=q�$  u&PH�=��$ 1Ҿr�B 1���{��H�R�$ H�K�$ Z�H�B�$ �S��H�� H�=*�$  u,H�=y�$ 1�H����H��H��H�zH�= �$ ����H���$ ��H��{�B �    1��^���I�ຉ�B 1�H�-�$ H�5��$ H�=��$ ��|��H���$ H�� [�ATI��US1�H����H��A�|�@��t��������1����������W�H��H�l$$�2�����B �   H���1��e|���;H������H9�u��=8% 1������=>�$ �����=&% �����<��9f H���}���H��u��=N+% �k����A+% ���]����=2+% �Q���H��[]A\�ATUS�   H�� �j�����u�H�\$L�d$ H���T���H�ÈC�L9�u�W�$�=1�����B �   H���1��{��H��H������1҅�uq����1����^% �������d�$ ��������J% ����������9f H��H��u������������������������   ���ÉM*% H�� ��[]A\�P����Z<����ÿ   �L���AVI���������AUATA��9f US1�A�<$ �c  �+������;f 1��y������;f �n������;f ��������;f ��������;f �8������;f �,������;f ��������;f ��������;f ������ <f ������<f ������<f �������<f �������<f �������<f ��������<f H�������H��u�1틼�0<f H������H��u닻H<f 1��������L<f H������H��u닻\<f 1��~�����`<f �s������d<f H���d���H��	u�1틼��<f H���M���H��u�1틼��<f H���6���H��u닻�<f H���;f A�   �������<f �������<f �������<f ��������<f ��������<f ��������<f ��������<f ��������<f ��������<f �������<f �������<f �������<f �������<f ����H��  H��tH�� �d H��I���1��e�����  H���V�����  �K�����  �@���A��tA�   몋� =f �(���H��H  I��H��   �z���[]A\A]A^�AUATA��9f US1�RA�<$ ��  �X���1�����H�H���;f �������;f �������;f �������;f �����f���;f ��������;f �k������;f �`������;f �������;f ������ <f ������<f ������<f ������<f ������<f �|�����<f �q������<f H��H��u�1��Z������0<f H��H��u��E���1퉃H<f �8������L<f H��H��u��#���1퉃\<f ������`<f �������d<f H��H��	u�1����������<f H��H��u�1����������<f H��H��u������H���;f A�   ���<f �������<f �������<f �������<f �������<f �������<f �y������<f �n���H�H���<f �`������<f �U������<f �J���H�H���<f �<������<f �1������<f �&������<f ����1҅�~H�Hk�(H�� �d H��  H���������   �������  �������  A��tA�   ������Hǃ�;f     �� =f Hǃ�<f     Hǃ�<f     H��H  I��H��   �Z���X[]A\A]�AUATU1�SRH��% 9-�% ~H�;��H���������{������{�������{�������{�������{�������{�������H�-C% E1�D9%1% ~v�}E1������}�����}����J�\-f���t9Hk�H�% �;�������{�}����{�t����{
�k����{�b���I��I��u�A��H��X�X[]A\A]�AUATU1�SRH��% 9-�% ~[�]�����H�����C��L������C��A���f�C��8���f�C��/���f�C��&���f�C�����H�C�    f�C�H�C�    �H�-?% E1�D9%-% ~{�����E1�f�E�����f�E�����f�EJ�\-f���t;Hk�H�% ��������������C����f�C����f�C
����f�CI��I��u�A��H��X�|���X[]A\A]�UH���������SRH��"% H��`if ��  H�{"A ��  �   ��������H���7����{�����{������{ ������{(������{0������{8������{<������{@������{H������{P�����{X�����{`�����{d�����{h�����{l�����{p�����{t�����{x�z����{|�r������   �g������   �\������   �Q���H���   H�� �d H��H���6������   �+������   � ������   �������   �
������   ��������   ��������   �����H���   1�H��tH-�;f H��i�����x��������   �������   �������   �������   �������   �v������   �j������   �q���H�[�,���X1�[]�����SH�=� % H��`if tH�_H�"A u�"�������  H�����h-  ��������N  <�2  ����1Ҿ   ��   �L�  H��H�������'����C�����C�����C ����H�H�C(����H�H�C0������C8������C<������C@�����H�H�CH�����H�H�CP�����H�H�CX������C`�����Cd�����Ch�����Cl�����Cp�����Ct�����Cx�����C|�������   �u���H�H���   �g������   �\���H�Hk�(H �d H���   �D������   �9������   �.������   �#������   ����H�H���   �
������   ��������   �������~"��H�Hi�H  H���;f H���   H���;f �Hǃ�       �������   ����f���   ����f���   ����f���   �w���f���   �k���f���   �w���H��Hǃ�       Hǃ�       �|������   H��Hk�\H�jd H���   H�CXH� ��@H�C"A �S`�Cd�=+  �����𿭵B 1��:>������[�SH�T% H��`if �.  H�CH��uH9� Gf �"  H��H��u��   H=C�@ �  H=)�@ uM�   ��������H�������{�_���H�{ H+=�% H���K����{(�C����{,�;����{0�3����\H=��@ ud�   ��������H���?����{�
����{����H�{ H+=% H��������{(������{,������{0������{4������{8�.  H=�-A u{�   �O����S���H�������H�{H+=#% H�������{ �����{$�����{(�z����{,�r����{0�j����{4�b����{8�Z����{<�R����{@�J����{D�   �   H=��@ tH=0�@ uP�   ���������H���C���H�{H+=�% H�������{ ������{$������{(������{,������{0�FH=[�@ uC�   �g����k���H�������H�{H+=;% H�������{ �����{$�����{(����H�[������   [����1���������H��������S�2���<��  ���$�еB ����1Ҿ   �H   ��  H��H��������c����C�[���H�H��H�% H�C �E����C(�=����C,�5����C0�-����C4�%����C8�����C<����H�{ �C@H�C H�XhtH�CC�@ H���(  H����l���F�������1Ҿ   �@   ���  H��H���%���������C����H�H��H�% H�C �����C(�����C,�����C0�����C4�����C8H�C H�XhH�C)�@ �d  ����1Ҿ   �@   �i�  H��H�������D����C�<����C�4���H�H��Hv% H�C �����C(�����C,�����f�C0�����C4������C8H�C H�XhH�C��@ ��  ����1Ҿ   �H   ���  H��H���$�������H�H��H% H�C�����C �����C$�����C(�����C,�����C0�����C4�y����C8�q����C<�i����C@�a���H�{ �CDH�CH�XhtH�C�-A H���\&  H���k��������d���1Ҿ   �8   �1�  H��H���q�������H�H��HN% H�C������C ������C$������C(������C,�����H�C��@ �C0��   �����1Ҿ   �8   ���  H��H����������H�H��H�% H�C�����C �����C$�z����C(�r����C,�j���H�C0�@ �C0�W����1Ҿ   �0   �\�  H��H�������7���H�H��Hy% H�C�!����C �����C$����H�C[�@ �C(H���%  �Y����𿙵B 1��8���E���[�S����  1Ҿ   H�H���<�    �% ���  �   ��H��% �l�  H�5y% �=�% 1�9�~�������L����L�H�����[���  �=��$  uH� �e �    P1�H�׾ �e �   �1��":���   �$�e �   �:��� �e ���$    Zø �e �AUE1�ATU��SR�?�  �   1Ҿ   H�H��1�k�8�b% ���  HcV% �   H��H�;% 1�Hk�8H������  H�"% I��D9-$% ��   H�{% I�$I�L$H�5q% H��H�I�T$H��H��H�CA�D$���CA�D$
���CI�D$Hk�XHx% H�LHH�C Hk�H�H�KH�IH�K(�@t/��H��H�TP��x9n% �����	Hk�H�DH�C0�H�C0    A��H��8I���/���X��[]A\A]�S�  S����  1Ҿ   Hc�H���=�% �����  �   ��H��% �e�  Hcn% H�=�% 1�H��1�H���1�H��% �=K% 9�~fD���fD�D�fD�DfD�D�
H���݉�[���  AUE1�ATA��USR�o�  �   1Ҿ   H�H��1҉ǉ% ���-�  Hcp% �   H��H�Q% 1�H��H���D����  H�-7% H�XD9-<% ~Z�C�H��A��H�����E��C����E��c6  H�{H��f�E��R6  f�E�f�C�f�E�f�C�f�E�f�C�H�E�    f�E��XD��[]A\A]���  S����  �   1Ҿ   H�H��1�k�4�}% �^�  �   ��H��% ���  H�v% D�W% 1�A9�~r����
�H���J�H���J�H���Jf�Hf�J01��|���|JH��H��u�f�Hf�J21��|���|J H��H��u���H��4H��뉉�[�!�  AU�   ATE1�U��SH���Q�  ��H����  �
   1�H�H��I��E9�}`�=L	# f�St�J�f��w�   H�੿ u;f�H�|$A��H��
f�D$f�C�f�D$f�C�f�T$f�D$
f�C�f�D$�8���뛉���  H��[]A\A]�AWAVAUE1�ATA��USR��  �   1Ҿ   H�H��1�k�X��	% ���  Hc�	% �   H��H��	% 1�Hk�XH���D���a�  H��	% H��D9-�	% �	  f�Ef�Cf�Ef�Cf�Ef�CH�?	% H�U L�<�H�UL�;L�4�A�6A+7L�s�sA�~A+�{��u	�C4   �&��u	�C4    ���B����~	�C4   ��C4   A�A�9�}�C,�S0��S,�C0A�GA�V9�}�C(�S$��S(�C$H�U
1�f�SH�Ef�C f���tHk�H�% H�JH�K81�f���tHk�Hu% H�PH�S@A��H��H��X�����XD��[]A\A]A^A_���  AUE1�ATU��SR��  �   1Ҿ   H�H��1�k���% �N�  Hc�% �   H��H�% 1�Hk�H�������  L�%�% H�XD9-V% ~f�C�H��A��I����A�D$��C���A�D$��3  H�{fA�D$��3  H�{H��fA�D$���2  fA�D$�H�C�H��H�% I�D$��X��[]A\A]��  S����  1Ҿ   ����  ��H��H�N% ��  H�B% �   H�PH��% ����v% �P���e% H�PH�@H�Ӊz% 1��؉�% ������  Hc�H��H�t% 1�H���[�AU1�ATUSH��H�0% �5�% H�=;% 9�~H�H
��H��Hk�8H�LH�IH�H����;�$     1�1�1�H��% D��% A9�~)H�z8H�J@�GpH��tH9�u����Ap����H��X��҄�t��$ ��$ 1Ҿ   �<�    �X�  H��% �5�% 1�H�Sp9�~Hc:H�B��H���B�    H����=+% 1�9�~OHk�XH"% H�H8H��tLcIpL�AxL��K���QpH�P@H��tH9�tLcJpL�BxL��K�����JpH���1�9-% ��   H��E1���3��D9cp~/H�CxH��N�,�I��I�E �P�0��3��I�EH��P�0��3���ˋ|$�L$A�   ��A���CHD�$�t$A�0�A���CL�k% A)�A��    D��% ��A9�A�@�)։C �    ��    ��H��s$�3% �5Q% )׍�    ��9��F�)щC,�    ��    ��H���H�뀉K�����H��[]A\A]�AU�-   ��ATH��"US��H��8H���$ 1����$     ���$     ���$     ǀ�<f     HH  ǀx;f     ǀp;f     H=   u�Hc��$ �L$Hi�H  ǀ�;f    �Z�  �   �   �>�  �  �=�# �L$u"��B ��	~��B �	   H�|$1��X������0��0�D$E�\$�D$M�L$�D$ H�|$���  ��%     �ōx
�#����}D�e	�����}�K����}�%����}�����}�����}�����}�T����w�����% D����  ��Lc����D9��   D����  H��% �   ��`f �߾   D)��4�  D��H��H��% �j�  ���$ L-% 1��D$,J ��   �D$ �   H��!H�D$$L��։���H�������t� ����@�p�9�v��vۃ�~<H�=x6$ �   ��1���B �e����V�B �0���K����I��%  L��������$     �}H�s% �_f �����=O�$  t.1ۃ<��9f  tHi�H  ��Hǀ�;f     �}��H��H��u���$     � %     �  �=�#  t�`-  H��8[]A\A]�P�A  �.  �@3e Z�[  �J��u�   ;:tW�B ���"�BD�B��u�   D9�t9D9�����Å��������+:D)���������1���9��������AUI��ATUSH��AP�w�{����:���{A�u������:��)�t8�s�;A+} ����:���sA�}+{A������:��Y��[A�<]A\A]��:��Z1�[]A\A]�AWAVAUATUSHc�H��(�� % 9��޿j�B 1��*��H��H % D�sH�[
Hk�8H% E���r  L�K ��$ A9AHu	H��8A����A�AHI���`f M�Y�hD� ��D��������`f E�SE�A��D��D������A9�t��5� % A)�E)�l$�=� % H�T$D�T$D�d$D�\$�L����5� % �=� % H�T$A���3���A9��g���I�y@ u1���   A�At�L�{0L�c(I�I9$�=���A�oE�/A9l$ANl$E9,$EM,$D9�~�H�t$��`f �9�����A�A9$t&��D��+=" % �T$�E9��9? % �T$}�3 % A�GA9D$t���+=��$ �9��9 % ~���$ � % 9��$ ������>����   H��([]A\A]A^A_���s���u1������������USPHcߋ5��$ �=��$ Hk�4H5�$ H�������Ń�u1�Hc��|C0������tE�5y�$ �=w�$ H�������9�t(��Hc��|k0��s����u1�������Y[]�t����   Z[]�H�GXH���$ ���$ H� H)�H����H�FXH� H)�H���$ H��Љ���Hc����r|�Wl�G �Nl���$ ����7$ D�G)ЋV ���$ �)�D���$ )��F���$ ���$ �O���$ �V)ȉ��$ ���$ ��$ ���$ D)x��j�$ �����w�$ 1��AUATUS��[e RH�m�$  af ������   H�kL�cH���t1�l(  ����   L�-?�$ L���(  H��A�EL�-)�$ �(  �+�ƽ  ��tjL�-�$ L����'  H��A�EL�-��$ ��'  A�EH���$ ���B+B���B��L��H��B 1��&&��H���$ �SH���P�H���$ H���9���X[]A\A]�Hc�Hc�Hc�H��H=
�$ H�GxH��H�DPHk�H��$ �Hc�Hc�Hc�H��H=��$ H�GxH��H�DPHk�HS�$ H�@�Hc�Hc�H��H=��$ H�GxH���@����1��GtH�G8H9�uH�G@ËD�OpI��1�A9�~!I�@xL��H�<������H��t� 9�O�H���ډ��D�OpI��1ɺ  �A9�~!I�@xL��H�<�����H��t� 9�L�H���ډ��AWA��AVAUI��ATE1�U��S1�H��hE9ep~KI�ExL��J�<��N���I��H��t.� D9�~'��t��u���B 1��$���A��A�Hc��ÉT�I��믅�t�l$1�H��9�~�T�9�O���H��h��[]A\A]A^A_�D�OpI��1ɺ���A9�~"I�@xL��H�<������H��t�@9�O�H���ى��D�OpI��1�1�A9�~"I�@xL��H�<�����H��t�@9�L�H���ى���Ƌ�$ H��$ Hc���9�~I��D�OH��I��fF9Lu������D�OpI����1�A9�~#I�@xL��H�<��%���H��t	�@9�O�H���؉��SH���   Hc�Hk�XHn�$ H��u[���   ��#w�� H��H���  f�Cf��Xt3f��
t+f��'t%f����  �f��at��  ��}f����  f�C��f=� ��  ���$�ظB �   ��   H���Y���z  1���   �U  �   �Z  1���   1Ҿ   �  1��G��   �@�   �H��输���0  1��  1Ҿ   ��   �   �  �   ��   �#   H���3�����   �   ��   �   ��   �   H���U���   �   �   �   [����1�1��wH��������   �	   �   H���V���   �   �t�   �mH���E����z�   ������   ������   H��� ����W�   ������   �/1Ҿ   H��������5[�5���H���F  H����  ��
   H���_}����   H����T��f�C  �  �   ��   H��[��T��H��[��U���   ��   H��[��W���   �Ҿ#   �1�H��[�������   ��   �   1��   �   �   �   �1�1��n1Ҿ   �eH��[����1�뙾   �t�   �m�   �f�	   �_1Ҿ   �3�   �O�   �H�   �\����   �R����   �H���1Ҿ   H��[����H��uH��[�  �   ��
   H��[�0|��[�SH���    H��f�Fuf��.t#�Of��.tf��/t)f��u=�   H����{���#�   H���V���   �1Ҿ   H������1�H��[�  [�SH��H�?H�GXH��9G ��   �r�F�f����   ���$�8�B ���$ �
   ��CD��   ����$ ��CDu}�   1�1�[�^����{D u�t�$ u_�   1�1�H�;���P����~��E���   f�B  �7���   ��<�$ u�   1�1��	����{,
[�������B 1�[���[Ã=:�$ ATUSu���$ u�p���L���$ L�A% � af L�A% I9�v?HcqD�A�yA�89�~&���$ ��y���D9 tA���A��H����H����5*�$ H�+�$ 1�9�~$H�Šcf f�z0uH�RHk��   H���ػ�ef ��gf E1�C����   �ȉCu~�C��tA��t!��uRH�H�P�CHk�H��$ f�B
�6H��SH�@Hk�H��$ f�P�H�H�P�CHk�H��$ f�BH�{�   ��  �   H��D���H�� H9��c���[]A\�AWE1�AVAUATA���USH��H�|$H�|$D������A�ą���  Ic�H��H��$ H�{h u�H�CxH��H�8�����I��H��t�Hp1��0H�5�'$ �*�B ����A�   �  I�VxH��H��H�R@H9�u	9���i  H����   H�5�'$ ���B �ʡ���=C�#  ��   �   ���B �)�#     �+�$     ��$    �E!����~hH���$ H����e H��H�<�H�,�    �gH��H�k�$ ���e H�|(�QH���N>% 9Б$ |"H�=�&$ �   ��B 1��������$    D�=��$ D�-��$ �D�:D�j1Ҿ   �@   ��  H��H����  I�nh1Ҿ   H�E��@ �@   H�E   L�u �E8 �  fD�m0H�E(   D�}4趷  H��H���  H�khH�E��@ H�E    �E(����H�] �E8 �  D�}4A�   ����H��D��[]A\A]A^A_�USR�5�$ ��~!�=:�$  t���$    i�4  ���$ �
���$     H�_�$ 1�9-g�$ ��   f�Cf����   ��f����   ���$Š�B H���9����o1��P1Ҿ#   H��舋���Z1Ҿ   H���w���f�C �CH�������9���$ �1H���U���'�   뷺   �   밉�H����U���H���t�����H���M���f�)�$   1�9i�$ ~QHk�XH�d�$ f�|(0u9f�=�$ ?~���B 1��M��H���$ H-7�$ H��H�,ՠcf ��f���$ H���1�H�� Gf     H��H��u�1�H��@^f     H��H��u뺠ef 1�H�׹   H�� �H���gf u�X[]�AUATA�   USR�w�" �����tE1��A��G�d$�`^e 1��Ef��u ��Hc����gf ���������$ X[]A\A]�D9�-H��D�k�|  Hc�H�}	Mc���gf ���c  B���gf H���1����ef  t	H9��ef tiH�� H=   u�E1�M��Ic�I��A���ef  u1H��L���ef H���ef ���ef ���ef ���ef H�G8H��0I�@�I��I��u��(�B 1������ATA��UH��S��uf�G  H�E1�Hk�HO�$ f�}�xD�@@��D�H
���$ ��� 1�Hc�9���   ���gf 9�uKH�=��$ �  ��H�E��Hc�Hk�H��$ ���gf f�PE����   ���gf �#   1��   D9�uGH�=��$ �1  ��H�E��Hc�Hk�H��$ ���gf f�PE��tp���gf �#   �   �QH��D9��G���H�=2�$ ��~  ��H�E��Hc�Hk�HM�$ ���gf f�P
E��t���gf �#   �   [H��]A\�-���[]A\Å�t1�f�~|��  H���    u.1��F ��  f�Vf��"�z  H�      H���f  f�F��f=� �P  ��SH��H���$�P�B H��H���O���(  1�H���&v�����  1��  H���.�����1�H��������H�����  �    ��   �   H���Ӹ��븾   �1Ҿ   ��1Ҿ   �ݾ   H���ar���1��d1���   ��   H����I���o����   �@1�H������������r  �	   볾   �1�먾   ��   ��   ��   H���L������1Ҿ   �M����   ������
   �a����   H����M��������   �E����   H���SL������   ��   1�H���#I����1��   �   �   �   �Ǻ   �   �a1�뷾   �h�   ��    �   �C�	   �N1Ҿ   �3�   �>�   �7�   �u����   �k����   �a���1Ҿ   H���E����U����
   H����p���C����   H����L���1�����   ��#   H��襆���   H�������   [ø   �����   u6��t2D�GH�5��$ 1��=��$ L���$ �H��H��fD;Dt
H��9��1��AVAUATUSL��H��`if �#  H�}"A ��   ���   )��   H�MXH�	H)�H��H9���   H��D�bD�jD�r �uH�ߋU�e�����u1���   �=��" t�C`�C H���   H��t	�P S �P�'   D��D��D���%����#   H����z  �E8H��$ �S ��k<��'   }k4���B u�����#   H���z  H���    t
ǃ�      �E8H�Cp    �Cx    �C8�   �(H�m�����H��H��fD;D�����H��9���$���[]A\A]A^�H�F�$ `if H�3�$ `if �H�+�$ H�xH�H�G`if H�=�$ �H�G������SH�
�$ H��`if t2H�CH���uH�SH�H��H�H�P���  �
H��tH����H�[��[Ã="�$  un�=Y�$  St%�,�$ �$ uHc��$ Hi�H  ���;f u=1ۃ<��9f  tHi�H  H���;f �  H��H��u��V����:���诫���@�$ [����H�[$ ATA��UH����S��4��"��H�U �4���B D��Bp�q"��H�U Bt[]A\�USH��RH��xp���R"����H��xt���C"���   ���=   OC(���   u	�=��$  uH��C B �C�   i��$ �  �   ���  �4���B �������!���{ uQ�K$�S ʁ�  ) ~
H�C   ) ���� ~�S ��C  � ���C$   �S$��t�� @  �   DщS$H��S Q ЋQd�C�� ��9�|	��   �SX[]�SH�H���w�H`��p89H �p8���Љ��$ �W��t��t�������S��t �=��$  tH���H�ߋp8��   @�]���f�{ tH�;H���   h�d u��   [�v���[�SH���6����C =   ~-   �C �{ �� �C    H��C$    H�ߋH`9H �����T�$ �,���H���   H��tLH�;H9�tD�w�H�P��"  H��ƋQ8)֍��q���:���v�A8����q����8���HЉQ8����   ��t�ȉ��   �Ct�C   [�H����   ����������   D����   ��t$�Gd   ���   �u�����S���   H����t
�ȉ��   ��V���H���O���H�H�@XH� f�x tH���F����{ y�C �K��tu��������u!1����    t�C|��u	�{< E���   ���" ��u��u���    t�{|�   EƉƃ���    t9C|t�p���w��t���   ��t���    uH���]���ǃ�      �
ǃ�       H���?����C<��t���C<�C8��t�ȉC8�C@��t�ȉC@uH����   �����CL��t�ȉCL�CD��t�ȉCD���   ��t�ȉ��   ���   ��t�ȉ��   �C8��t=�   �tǃ      �(�CL��uǃ      �=�   �t�ǃ     [�H�$/% �jf �AT�G�A��U��S��if 9C}H�����39�~^��D9�~ND�����1  H���$ H�PH���$ H��H9�tH�J�H��H�J��H��H)�H��H��Hk��HЉ(D�`�k���1  �+H��D9c}Y�E�p��E�xD9��t1  H���ED9�|މC�D���[1  D�cH9�t!H��H9-�$ tH�EH��H���H�	�$ []A\�U���G�S��if Q9C}H�����39�~&��9�'�1  ��C�p��C�x9���0  H��9k|��
Z��[]��0  X[]����$ �����]% H���$   ����$ H��$ �if �UH��SVH�H�=�-% �p�8�3  ��H�E�p�8�#  A��A)���   �=�]% ��]% ��	( )��4�9�s)�A9���   �Ӎ)�9�r)����)�A9���   �ځ�   @��   @�����<�@�f �4�@�f 9�tmH�E0H�-% H��tSH���$ �9X~E�Y9}>H�H9u,H�������  H�XH!�H#QH9�uH��,% H�@f�x tY��[]�v���Z��[]����X[]Ë��% 1�9W}
1�;W�������% 1�9~
1�;O��������   H�ATH��UHc��ae Hc��ae S�,�Hc��ae Hc��ae �4�D�$��<���  D��+z\% ����  D�j\% �   D��)�A��A�xw�V\% �4�<9�s)�A��1�E9�v[���9�rD)Љ��)�1�A9�vC�ځ�   @��   @1�������@�f ��@�f 9�t�P���if 9P}H����1�9@��[��]A\þ   ���USHc�R���$ 9��޿��B 1���	��H��H��$ �c[% H��kH�[
�8H��$ Hk�8H��$ ;=��% }�P�p�%  H��d' �H��d'     H���$ �x;=R�% �p
95�( u�P��$  H��& �H��&     H�=��$ �>  �̓��tH��H��8�������X[]���s���u1������������USPHcߋ5��% �=��% Hk�4H�$ H����  ��H��|C0��Hc�����H�}H��H�������t�|k0��s����u1�������Y[]�Z[]�I��I��A��A�8@���t:A�H׍9y��1�A9�}D��)���~Hc�I�pI�:H���A�@M�D ��AW�   AVAUATUSHc�H��H�-*% L�4�H��)% H��H��)% �<����  H��H�*% L�$�H��)% L�,�1�A�F9���   A�|� �   �t�  M�L�A�    D�8C�E�~A9�DO�E��MI�E9�~IfC�<\ y<D��C�t] A�N
D�L$D)�A�T�H�$Hc�H�Hc|�H������D�L$H�$I���H���g���H��H��  ���B [�   ]A\A]A^A_�g�  AWHcǾ   E1�AVI��AUATUH�,�    SH��H�)% H��H��(% H��    H��(% �{��    H��(% L�$�H��(% L�,�H�T$财  H�KH��H�D$1�H����CD9�~qB�|� �   �6�  F�D��    �8E��B��{AI�9�O�Hc�D)�Hc�H��H��9�~&H�t$H��B�t� f�PfA�4L�rfA�tM H����I���E1��CH�|$D9�~eB�?��uH�޿��B �j����S<vEH��'% fC�|���   �(fC�D} �K
)�9�~D����B 1�����H�x'% �K
H�I���� �  H��[]A\A]A^A_�UHc�SQH��'% H�j'% #4�H��'% Hc�H��H��H��2�0��~�   ����  H��!H�'% H�<� u����H��&% H�H��Z[]�AW�   �0�B AVAUATU1�SH��H�D$? �S�  1Ҿ   D� H��H��B�<�    ��  H�D$A9�~-H�޺	   H�|$7H���m2��H�|$7�%�  H�L$��H���ο0�B �[�  �   �7�B ��  �7�B I�ċ �D$(肜  ��衜  �@�B �D$I�D$H�D$�͛  ��t+�   �@�B 蠝  �@�B H�ŋ�A�  ���`�  �D$��D$    1�1�\$(1Ҿ   �<�    �&% ��  1Ҿ   H�&% ��%% �<�    ��  1Ҿ   H��%% ��%% �<�    �ҟ  1Ҿ   H��%% ��%% �<�    貟  1Ҿ   H�f%% ��%% �<�    蒟  1Ҿ   H�>%% �t%% �<�    �r�  1Ҿ   H��%% �T%% �<�    �R�  ��WB H�P%% �:�  �I�B A���-�  �$%% A���%����u1��   E)��@   �[   E1�A�F>������C?����莇��D�sE9�|�    A���x�����]   E1���	�f���D9�|��   A���T�����H��$% ��H�D$��A�E
H��$% ����H��9�$% A���f  ��?u
�.   ����D9t$(uH�EI��H�D$�D$�D$H�D$D�0D9t$}�O�B 1��V��H�H$% Ic�L�<�    1�M�4�   L�I��H�D$ A�F��<�    ��  1�I��H�D$ I�UL�(fA�F�fA�EfA�F�fA�E
fA�F�fA�EI�F�I�E A�E9�~QfA�H�t$f�fA�Ff�BI�F���B��u!L��u�B 1��L$,H�T$ ����L$,H�T$ ��I��
H���I�}L�5�#% 1Ҿ   �M��U�  I�}1Ҿ   I�L=!#% ��8�  A�MI��   � 9��h�������H�|$�g�  �7�B 踚  H��t
�@�B 詚  1ۋ�"% 9�~�����������1ҍ<�   �   �Ϝ  1�H�#% �=�"% 9�~��H������1Ҿ   1�補  Hc�"% H��H��"% 1�H��H���9-w"% ~_H��"% H��    H�<�o�.�  1��5R"% H�w"% Hc�H��H�H��tH�P��H�K"% H��H�H�H�A    H� H��H��H[]A\A]A^A_�R���B ���  ��XB ���_"% ��  �   �ȉ"% +G"% �P�<�   ��!% 1��ʛ  1�H�"% 9�!% ~��H����X�U��WB S1�R虗  �I�B ����!% 臗  1Ҿ   �x��=|!% +=�!% �ǉ="!% ���h�  1Ҿ   H��!% �!% �<�    �H�  1Ҿ   H�$!% �� % �<�    �(�  H�� % 9� % ��~X��?u
�.   袃���=d!% �   �褗  H�!!% ������PH�� % �@����H�� % ����H���X[]�P���B 詖  �   ���R�  H�� % Z�P�g����.   �%����u����.   ����������.   ����Z�UH��SH��迕  ����uH�E H�t$���B �D$ H�D$1��P�����+� % H��[]�1��?-tLUH��SQ���  1��5 % H�) % Hc�H��H��t�   H��H���5�����u�C�	H�[�܃��Z[]��UH��SQ��������uH����B 1��������Z[]Ã=M�$  �o  AW�   AVAUATUSR�=�% 1�脙  Hcw% H��1�H���1�9��$ ~.H���$ H��H��H��H�L�H���$ H�T
����#%     1�9-#% ��~2�<+ t'=% �   Hc�Hk�(H -( �@�% 覕  H����H���@�  �=�% 1Ҿ   �٘  Hc�% H��1�H���1�9�$ ~<Hk�H�}�$ H��H�L�H�i�$ H�L�H�X�$ H�T
��Hc��' 1���5%     9-[% ~N�<+ uH����H�c% E1�L�,�A�ED9�~�KcD� �   I��H��Hk�(H,( �@�% �Ŕ  ��H���b�  �=��' 1Ҿ   ���  Hcv�' H��1�H���H�%�$ H=`if tH�x"A u�P<�H�@����%     1�9-4�' ~k�<+ uH����I��E1�I��H��*( L�D9(~�Mk�E1�LxC�|7=�% �   I��Hc�Hk�(HX+( �@'% ���  I��u�I���XH��[]A\A]A^A_釖  Ë�% �5�% S��)���   ���   ���nL% @����@�u��?  v���B 1�����Hcw% Hc@L% �5"I% H��+�L% Hc���f ��H�`�f �.% ��H�=7% �����H��@  ���H�=% ����������u�[Ë% �5% S��)���   ���   ����K% @����@�u��?  v���B 1��U�����K% Hc�% D�rH% � H��H��`�f +L% Hc�A����'.% Hc�Hc4���f Hc���f H�H�1҉�L�k% ��D�����A�<9L�L% A�<9@�<@�<H��@  ���u�[Ã=;%  Su
�.%    ��-% �P�;#% u	���% �% �5% ��)���   ���   ����J% @����@�u��?  v��B 1��W���Hc�% Hc�J% 1�Hc���f H�`�f Hc�n$ H�5Z% Hc�`be ���   ��=n$ �W��2D���H@  �hn$ ���u�[�USR�=_%  u
�S%    ��,% �P�;H% u	���=% �7% �5-% ��)���   ���   ����I% @����@Ǎ	u��?  v��B 1��y���Hc�Hc�% ��1�Hc�Hc���f H��`�f Hc���f H�H�Hc�m$ H�=m% Hc�`be ���   �Hc�m$ H�=J% Hc�`be ���   ��om$ �S��2D���H��@  H@  �Qm$ ���u�X[]ËN% �5D% S��)���   ���   ����H% @����@�u��?  v���B 1�����Hc% Hc�H% �5�E% H��+NI% Hc���f ��H�`�f e+% ��H�=�% �����H��@  Hc��H�=xH% �H�=�% ����������u�[�USR��% �5�% ��)���   �FH% ���   ��� �����u��?  v�ٿ��B 1������HcD% Hc��Ë5�D% Hc�Lc���f H��Hc<���f +}H% H��`�f ���*% I�H�1҉�L��% �����L��G% Hc�E�	G�
L��% G�
E�L��% A�	L��G% A�	L��% A�	�H��@  ���u�X[]�R�   1ҿ   ���  H�jG% �   ������H�XG% ��w1���r`@�� ���H�<G% �r@�� @�4H�+G% ��   ���   H�G% �H�
G% �� ���H��H=   u�X�R�5�C% ��C% ��C% ����9�@��@�u��?  ���   v�1�B 1��V����])% ��F% ��F% Hc=zC% ��
��Hc5iC% ��f1���	ЋpF% ����
f1�	�H��Hc<���f H<�`�f �50C% )Ή�A��H������A��Ё��  D	�L��(% A�L�+% A��O����u�X�R�5�B% ��B% ��B% ����9�@��@�u��?  ���   v�1�B 1��}�����(% ��E% ��E% �5�B% ��
��Lc�B% ��f1���
��	Ћ�E% f1���5oB% ����	ыiB% )�҉_B% Hc�Hc4���f J4�`�f ��A��L�d% H����A����ȁ��  D	�L��'% E�G�D�F�L��'% A�L�%% A��V����u�Xø@  1�)�����A% 9�~�����f H����1���@  t	��   )����~'% i�@  1�H�HY�$ 9�~H��`�f H��H@  ���USQH�=�h$ �=='% @  uH���N  �h�  H��h$     �9  H��u1Ҿ   � �  ��  H�xh$ �T�B �L�B �   �=��" HE���  L�Rh$ E1�M��@  E��I������A���  I�H��H��@�   L���L9�u�A��@L��@  A�� *  u�L��1��Zg  �   �]�B 訋  H��;p&% }�l&% �=�@% H��ߍp����2`  �ھ   �d�B 1��n�  H��96&% ~!�=N@% �5@&% H��5#&% ߃���_  �׾   �k�B 1��1�  H��9&% ~�5�%% �@% H��ލx����_  �ھ   �r�B 1����  H��9�%% ~!�5�%% �=�%% H��=�?% ރ��~_  �׾   �y�B 輊  ��%% H�q���?% �y��S_  �   ���B 蓊  �b%% �=X%% H��=o?% �q��'_  �   ���B �g�  �R?% �5D%% H��5'%% �y���^  �   ���B �;�  �5%% �= %% H��5�$% =?% ��^  Z[]�e  X[]�H�Qf$ H��tH���$ ��Hc�H�48H�H���Ë5�$% ��@  ��   ��   R+�$% 1��   ���A���@  )�Ei�@  ���E�A��D�������=�$% D��D�i�@  D)��v���E��@  A�   E)�E�D9T$% ~D��D���O���A��@  A���๨   �@  1�1�X��\  �9z~�z9z}�z9r~�r92}�2ËBD�B��uD����9:|lE���D�JE��uD9���Å������D1���+
D)�1�AT1�U��Sy
��D1����'D��H�Ӊ���� ���s
��A�������A9�����[]A\��H�H�RD�@���RD)�)�u����9�|a1������ATUS�Å�uA9�}�����;��D)�)ȉى�1�1�1�y1����$�׉������~����މ�A���r���A9�����[]A\�Ë��% A��A��1����% )�A)�A��E	���   AR��xmE��x2D9�~��D���6[  H�����B �   D��� [  Hcи���?�   )�9�~�����[  H�����B ���   ����Z  H�����B -   @�pD)ɉ�E��x1A9�}��D����Z  Hcи����FD���Z  H�����B    @�5)�9�~�Ή��Z  H�����B    �����|Z  Hcи����+���B Z�É=��% �׉5��% ����������% ��+5��% S��)Љ���1�)ȉ���1�)�9�|
9�t�ډÉЉމ������1�1�����[H�����B    @���4���B �����ø   @US��Q+�' �+?% ����=?% �4���B ������B ������>% �=B�' ������������  @ ��9�}$�Ɖ������   =   Mи  @ ��  @ OЉ�Z[]�Ë54$ �=f>% ATE1�U���S�K�����A��$��C ��   ~���?��  ��}
��=% ���-���
����5">% )Ɖ���  �����|ʋ�=% ��9�O�A��$@�f I��I�� @  u��5�=% 1���9�|%1ɉ�H��9<�<�f �����   @�� ug H����1틽��C ��������@�f ���uǅ@�f     ��B=% �H9�u��@�f H��H�� @  u����% []A\��=% �AUA�<   ATE1�US�   R�   ��  � ���.���D��������   )�����Oº    ��H���H�H�% I����4g H��H���   u�I��   A��I�� @  u�X[]A\A]���<%    �=�% �5�<% �USR���% ��<%     ��u�% @  �% �   �"��i��   �
   ����% ��������% �5�% A�   �=�% ��<% ��A���A���j<% A��D��;% A���{<% D���A��A��D�A<% A����|% A��D�<% D�B<% ��u9H�/�% ��A H�<% ��A H�1<% v�A H��;% h�A H��;% ��A �7H���% ��A H��;% ��A H��;% O�A H��;% #�A H��;% ��A �F��������>;% �@  ���������( �  @�����% �/�' 1�9�~f�� ��i H����1۽   ��% �=�:% 9�~<��ދL;% ��)����� �  ����1�)Ɖ����������������� �h H���1ۋ�:% 9�~4�� ug H���# �   �����4���1�)������� �g H����:% 1�A�<   1�L�>% A�   A�   ����1�i�@  ����A��D��)���AOÅ�H���H�L�H����g H��H��0u�H�ǀ  A��H��   u�X[]�P������.   �m���.   �m���.   �m����# �:%    �A�% �\$ �!:% �  �.   ��l�������.   ��l���-  �����.   �l����9%     ZË!�$ ��uH�6�$ �AT�B�A��U��S��r$Hc�D���Hk�4H�$ H�������H��DC0�ր�[]H�A\H��H�$ �H�H�=h�% �B���% �B���% �l�% B8��   �i9% ���H9% �W�_�% ����B ��8% H���# ����8%     �(9% ��  ��t3H��' `g ��1�H�Hm	% H��% H��`g H��H��0u��H���%     ��8% ���# �P�;��������L�����  �  �v�����$ �x������c����  �Y����
"  Z�N����AWAVAUA��ATA��U��SH��9�|��x9�7% ~9=�% }D��D���B 1�����Mc��=x�% B9<���g tQB�4� �h B�<���g ������5�% �ǉ�B��@zg �����5<A' ��B����g �|7% ����B��`�g �B����g B��@zg �W7% B��`�g Lc��߉H7% B�4� �g �a���D�5�7% F4� ug ��H��# A���։T$B�<��6����T$D�=��% B�<���B w�% �։�% A������A)�H�i�% D�=�6% H��u���   ��HG�H���% H��D�-�3% �-�3% D�%�3% H��% H��[]A\A]A^A_�%�6% �z6% �@% S1�9�~f�� ��g fǄ ��i ��H������g 1���   �5�6% H��?'  �g H����6% H���% ��h ��   �H��# ���<��K����<���B �5J6% �l�% �3���[�؉�?' �AU1�A��ATA��U��S� �g Q95��' D�DD�H�{?' H9�vD9+uD9cu9ktPH�Ø  ��H= �h u���B 1��@���H�S�@  D�+H�@  ����H�CH�װ�D�c�k�H�?' �  ZH��[]A\A]�HcGA��9�A��HcƋOA��9�|A�ȉ�9�|LH���|�t�L��>' �@  A� �GA�@�GA�PI�PA�@I���  H��H��>' ��A�p��D�OD�GI��L���AW�G�AVA��AULc�ATA��UD��SHc�H���D$E��E9�~D9�|B�4� �g �T$D��I���y�����E�n���9�}A9��4� �g ��D��H���T�����Ic̉�A9�~9�|D�4� �g H����Lc�D9�}D9�F�4� �g I����H��[]A\A]A^A_�H�5J% AVAUH���jf ATUSH�� @  ~H�����B 1�����H�5�=' H�� �g H�� L ~H��C.+Jx�H�����B H��1��l���H�5&�% H���h H�� �  ~H����B 1��F���� �g E1�H9@=' �l  Hck;k�S  HcC;s�' ��   ��3% �m�' ���10% H�*% H�[% �=�' ��% �T+��+W  �L% �J% 9�.�5�3% �=�' �- 3% 4� ug �������H�% �D3% H��9k}��   H��% �-�% �   ,����z  H�|% �+<�% �1Љ[�% �C)R�% �   ���2% AHă�O�H�H��
H 5g H���% �CD�pIc��D�LckA�E�H��D�E9�|+B�L+B�t+D��B��+V  F��+W  I���W����Љ��z  H�Ø  ����[]A\A]A^�AUATU��SQH�H��% L�BL�R(H�+% L�J0L�I�HL���$ L�	% ��A�BH�Jf���D�a2% E9cu���	�	A9u����yH��' �g �$Hc�Hiɀ  H���g ���`3g HN�H���' H�G8�OH��' ��+G��G���' �Z�' H�G0���% H�( H�G(H�n( H�B �@tA�H�=�% Hc�A9AM��% ��A�BA9AANA)ȉ�% A�@�% H�o�% H��tH��% �5�0% A���Hc�0% 9���   H�S�' f�<B���   H�=/�%  �5��' u#��/   ����/HG�H���' H��H��% �=&% D�-�0% ����1҉�A)�D���5b�' HcC0% D�-�( �-% H���' �4P�(���H�x��  Hc0% H���' f�P����' ��/% �' �1���X[]A\A]�AVAUATU���SHc��' ;f�' ��  �b�' ���  �� ��i ��9�|�Y�=��'  �� ��g t'�s�D�A9�|�r�D9�|H�=��% D�D@��W  D�%�' A��A9�|D�b��=3�'  t%A�t$��9�|�q9�H�9' @�t��W  E1�=&�'  ts���' � ug �Ћ5��' D�-��' ���<���C �/������' �/   A)ŉ�A������/HG�H�`�' H��1�H���$ ���' ��.% �����+% �=��' ��tR���' D����$ D�%��$ �O% ����H���$ ��.% Hc6�' �@% fǄ ��g ��f�� ��i �I  �=3�' Hc�' ��to�B�' A����' �3�' �� ��g A��D9�D�r�D9�I���' D��:�$ D�57�$ ��% �����H��$ �K.% Hc��' fD�� ��i ��=��'  t
��f�� ��i �=��' �z�' ��tq�d�' ���  h�' �R�' Hc�������i 9�|�XA9�|K�n�' D����$ D�%��$ �(% �e���H���$ ��-% Hc�' f�� ��g ��=�'  tHc�A�D$f����g �=��'  tHc��' H���' fD�,P���' ���' ��' ���' ��' ���' ~�' ����[]A\A]A^�H�=�$ ��f �i  AWAVAUATA��US��H��9=�,% ~9�~D��޿?�B 1��N���H���$ H�AH�}�$ H�A f�H H���$ �A   @���' + �' �1�)к   @=   @O�)�H��Ջp�8�,�����Hc����ǉD$�4���B �U���H�d�$ ���' ���' H�A�$ �=�,% �XD�`<� ug H�A�D$�{�' �7���L�-�$ ���' A�ED9�};Icċ=K,% A)�<� ug �	���H���$ A�E�A+��' �A���F�' �A�A�EL�%��$ �5�% L�q�$ L���$ A�$E�\$�/�'     �)�'     A�z�'�'     ��D��)�)�f�|$���' H�d�$ ���' ��'     H�@8    M��uyL��H�=��$ B�<����'    ���'    �=��' H�=��$ �GtH�z�$ B���)�H����   �ARH�@(��i ���' H�@0@�i �@   H�p �*  A�8H�@0    H�@(    �@    9�~�@   �H �9�}H�   ���H�PA�PA9�}
�HD�X$�9�~�H�@$   �9�|�HH�@0@�i �@ ���A9��HH�@(��i �@$   �A��A��E�l$
A)�A)�D;- �' D�5��' D�|$D�=]�' uE�x
E9�uD�5��' A�   9�u!I���  ��  M�xM!�M#l$M9�A��E��D�-p�' D�-M�' A�   E9�u!I�  ����  M�HM!�M#|$M9�A��E��D�=b�' 9�}A9��#�'    �E�'    E9�}AM�BL� �$ G��D��' L�6�$ A�Ct	D�-��' �L���$ C�)���' 9�}-I�J
H���$ �����' H��$ �BDDl$D�-��' A�R��' ��' f�|$ tFH�#�% Hcd�' �j�'    H��H��H�H)�H�x8��' H�=%�' )�H�H�H�H���% �Z�' @�' .�' $�' �J�' ��   ���' ���' ��)�=   �v��)�=   @�   @�|$G����4���B �?�����' ���' ;��' x�؉��' H�2�$ H�5۶$ �B��' �Z(%    @)�H�=[�%  �M�' ueH���$ H�
H�R�@�rf���(% 9qu����291u����yH��' �g �$Hc�HiҀ  H���g ���`3g HN�H���' H�W�$ ���% 9|
��'     ;P|�@
;<�' t
�$�'     �5��' �=��' �=��' ���5��' �1���D�%`'% �5��' �=��' ��A�����' �����5Q�' �=�' A)�D�%a�' �����D�%!'% �5��' �=)�' ��A���i�' �����A)�H�=��$  D�%"�' ��   �=6�' �=��' ��;=*�' �= �' }9D�%�&% �5Q�' ����A���5�' �=��' A)�D�%:�' �g����؉��' �=��' ;=��' ~9D�%�&% �5
�' �?���A���5��' �=��' A)�D�%��' � ����؉��' �=��'  t"�k�' �5��' H�="�% �P��w���H��% �=��'  t"�@�' �5f�' H�=w/' �P��L���H�h/' ����H���$ �B��H�' tXH�z( uQ���' H�D- H�=��% H����i )��Hc��H���% H��H)�H�q�$ H�H(���' )�H�H�H�H���% H�O�$ �B����' ��   H�z0 uO���' H�H�=f�% H����g )��Hc��H�O�% H��$ H��H)�H�H0�T�' )�H�H�H�H�'�% �=x�'  t1H���$ �P��u���@$   ��P�P��u���@ ����PH���$ @H��[]A\A]A^A_���[�'   d �AWAVA��AUA��ATA��U��SAP��w��vD��_�B 1������;-\�' ~�-T�' ��Hk����i E��un��uH�50�' �UA���B ����Hk����i uH�5�' �UA���B 1�����Hk�D+%��$ 1�ǃ�i     fD��C�i D����i H��H��u��y��uH�5��' �UA���B �4���Hk�E�~�ǀ�i    Hk�L�f�� �i �tH�5��' A�N0�UA1���B �����Hk�D+%4�$ Hk�L�fD�� �i E����i X[]A\A]A^A_�H��H�8 tH����H)�H����' ���5  AW1Ҿ   AVAUATUH����S��1�H��(�fm  Lc5��$ H�� ( �P�$ M���D$Ik�(H�D$9��' ��  H�D� ��i �,  E��H��L�l$���' ����H���' ���D9d$��   L�5� ( H�5��' �   M�L���(U����ugA�vA�VD����A��0�=�t$  tL���T$�t$�h  �T$�t$��1�����H�� ( L��p@��t�P��A�   D���0����A��I��(�`�����' I��I�����uH���' B�     ��   ��E1�E1���' �=��' D9�~zA���i ���t��u^A�EAE1ɉD$�"H�5��' A�UA�K�B 1������8I��I��t/fC��N�i �u�T$�{�B 1�L�L$H�5`�' �����L�L$��A��I���{���L�-��' �   1�M�A�} k��k  Hc,�' ��i I�EH���' Hk�J�D H���H���"���H��([]A\A]A^A_��1�fǄ @�i ��H��H=@  u�����H��' ��i �H��' H=��i tH�PPH���' ø��i �USH��R�-!% �<���   �h�' �s��������' ����  �|2�Hc- % H�5�' �����J�$ H҉=E�$ �49�|�Ή55�$ H�5B�' �9���$ ��$ 9�$ ����H�S)�H���$ �=�% � % �CH�\�O����-j% X[]�AU�   ATUSH��R�=��$ {8��f  H��H�C@H���$ H��uH� % H��% �6�CH�   t,H��% ��%   H��% H�W% H�� ���H�(% �S0�C0��% �{4���s,D�-|% 1Љ=�% D�c()Љ5�' ����% �%���A)ŋCD�-v�' ��% ��% 9C|:E��A��x	�E D9����B 1��n���Mc�Jc|�H��:�����% Dc0�H��% H��% X[]A\A]�AWI��AVAUATUSH���_�5�% +�% D�o��D+-�% �����5�% D��A���t���A�A���� �@  �=�% D��A���d����5R% �߉��C����5�% D����3���)É�����1�)�D9���  A�w<;5�' r���B 1�����E�o<A�W@L���I��L-��' %�  A;E |��B 1��[���E�g@A���  Mk�MeA�<$ t'A�wA��L���A+G8-   p��E�tDA�D�E�t$A�D$�D$H���$ Mc��B+����n����% A��A��D9%,% �0  H���$ ��B�<���@���X% �������	  �h����\% H�a�$ H��A���   �CH�����C,A�G�CA�G�CA�G �C B��C$+C�% E��C4�    AIĉC��% 9��p��s�   ��������|$ tH�G�$ ��B���ʉS(��C(    �C0�CD9�~
D)��C0C(D�s8A���   t
H�C@    �DH�ǻ% H��u4H��$ A�GA�u&�   +}% �/   ����/O�H���' Hc�H��H�C@H��[]A\A]A^A_Ë}�# 9GXt^S�GX�Gf���6% yH���' �g �$Hc�HiҀ  H���g ���`3g HN�H���' H�_`H��tH�������H�[(��[��AWAVAUI��ATUSH��XH��0;5}�' r���B 1�����I�E ��PH�މ�H��H&�' %�  ;|��B 1������I�E �5�' �@%�  Hk�HCL�pD�`A�EL����  `�H�r�$ B+�������)% A��A��D9=�% �!  H���$ �5 �' B�<��������% ��������   H��$ A�M�    �D$H    B+�� �d )�E���D$4AI��j% �t$9��P���% ���' �T$���D$,�[�' E��t�؉D$0H���$ B���ȉD$(��D$0�D$(    D9�~��D)��D$0D$(H�[t% �l$8�@@=�   �tH�D$@    �2H�o�% H��u!I�E �@�t	H���$ �H���' H��x  H�D$@H�������H��X[]A\A]A^A_�SH��s% H�H�@XH� �@f����% yH�`�' �g �$Hc�HiҀ  H���g ���`3g HN�H�:�' H��   H��' ��i H�l�' @�i tH��  ����H��(   tH��(  [����[�H�~�' H�t$�H���������H��H����i H��H�ȸ��i A�Ʌ�u�H9�vH��PH��`���H�@�H�H���H�5��' H��P1�H�D$���i H�rH�T$�H��'  �i H��'  �i D9�}`H�D$�����H��H9�tD�B,A9�}D��H��H�R��H�8H�P��H�:H�8H�WH���' H�@ �i H�H���' H���' H�B��AUATI��USR�WHcG9�|fǄ ��e ��fǄ @f ��H����H��$ H�h�A�T$A�t$H���jf �\  �]9��H  D�mA9��;  �} uH�}8 �*  9�EL�A9�DO�U9��щ�A�L$,9�~H�}8 ��   D���H���X�����   9�~A�t$A�|$H�U ������tȋE�} A9|$ |����M$A9L$$�������   ���u,Hc�A9���   f��6@f �uH�E0f�pf��6@f H����Hc��u%A9�|hf��6��e �uH�E(f�pf��6��e H����Hc��u@A9�|;f��6@f �uH�E0f�pf��6@f f��6��e �uH�E(f�pf��6��e H����H��@�����1�$ Hc�9�|-f�� @f �uf�� @f f�� ��e �u
fǄ ��e ��H����H�
�' @f L��H�\�' ��e X[]A\A]�b���S����H�=�' ��i wH�&�$ H�X��7H���' H�� �i t�H������H�[��H�{8 t�S�sH������H��@H���jf sރ=�%  u[����[�AWH�V@AVAUATUSH���H�|$��D$ȋG�D$ЋG�D$ċG�D$̋G�D$�H�D$؊H��H���H��N��H��N��H��N��H�H9�u�D�T$؋D$�D�D$�D�\$�A���y�Z�D$ȋ\$�A���t$ċl$���D��D�d$�D�l$�ЋT$�3T$�A���y�Z#T$�3T$�D$ċ\$�D�t$�D�|$�D1�#D$�3D$�ȉэ�3�y�ZD�L$���ȋL$���1�!���D1�F���y�Z��������1�!���1�A���y�ZD�A��A��D�A��A1�A!�A1�A���y�ZAȉ�����Aȉ�1�!���1�A���y�Z�D����щ�1�D!�A��1�A��?�y�ZD�|$�����D1�!���1�A��7�y�Z������D��1�!���D1�G���y�ZD�$��������1�!���1�A��	�y�ZD�L$D�A��A��D�A��A1�A!���A1�A���y�ZD�L$Aȉ���Aȉ�1�!���1�A���y�ZD�L$�D����щ�1�D!�A��1�A��9�y�ZD�L$����D1�!�1�A��1�y�ZD�L$��������D��A1�1�E1�D3T$A1�!���D1�G���y�ZA����������1�!���1�D�D�A��A��D�A��A1�A��A!�A��A1���E�D�L$�B���y�ZA��E1�A1�D3L$A��A��A!�A��D1�A1�D���E�B���y�ZD�$A��A1�D3D$A��A��D�D$�A���\$�A1�A!����A1�E�A��B�� �y�ZA��A1�E1�D3D$A!Ӊ���E1�A1���A��A�D�B���y�ZD��A��D1�3|$��D1���A1���A1����A��F�����n�t$�1�E��1���D1�3t$3t$�A����D��D��)���nD���D1�3L$1�E��D1�D1�A����D�A���D��*���n�T$��3T$�3T$D1�E��1�D1���A��D��A��E�ލ�(���n�$E1�E1�A��D1�A��D1�A��1�E����B��3���nD�t$�D3t$E1�A��A1�A��A��D�t$�E��E1�A1���E�D�|$�E�G��3���nD�4$D3t$D3t$�E��A1�A��A��D�t$�E��A1�A1�E�D�|$�E���G��5���nD�t$D3t$E1�E��A1�A��A��D�t$�A��A1�E1�A��E�D�|$�E�G��4���nD�t$D3t$A1�D3t$�E��A��A��D�t$�A��E1�E1�A��E�D�|$�D�B��5���nD�t$D3t$A1�D3t$�A��A��A��D�t$�E��E1�E1�A��E�D�|$�D�B��3���nD�t$A��E1�A��D3T$�A1�D3t$�A1�D3T$�A��A��D�t$�E��E1�D�T$�A1���E�D�|$�A��E�G��3���nD�t$E��E1�A��E1�D3L$�A1�D3t$�A��D�t$�E��A1�A1���E�D�|$�A1�E1�A��E�D�|$�G��5���nE��E�A��E�D3L$�A1�D3D$�A��G�����nD3D$�D�L$�A��D�|$�E��A��E1�A��E1�D�A��E�F�����n�l$�E��1�3l$�3l$�A����1�3|$�3|$��l$�D��D�|$���D1�D1�D�A��D�E��E�荜+���nE1�E��E1�A����A��D��G�����nD1�1�1�3t$�E��1���A��D1�3L$�D���F�\- D1�A��A��;���nD����1�A��E�L$�D1�A����D�|$�D�A��3T$�3T$�A��2���nD1�1�E�A��1���D�t$�A�����T$�D��D�1�D�\$�D�T$�A��	���n1�A��A��D�3D$�3D$���D1�E�D3t$�D3t$���A�����nE1މÉ�A��	�A�!�A������!�D	�A��A��D�A�� ܼ�D�D$�D3D$�D�t$�D3D$�E1�E��A��A	�A��E��A��D���A!�A!�E	�A��A��E�B��ܼ�A��A	�E��A��A!�A!�D���E	�A��D�t$�D3t$�A��E1�E�A1�B��ܼ�A��A��A	�D�D�t$�D�t$�E��A����D3t$�A!�A!�A1�E	�A��E1�A��A��E�D�D�t$�B��ܼ�A��A	�E��A����A!�A!�E	�A��A��E�F��ܼ��T$�3T$�D1�3T$��T$���D�\$�	�!�D�A�щ���!�D	�E��A��D�A�ɋL$�3L$���ܼ�D��3L$�3L$�D	���!��L$���D��A��D!�	ȉ���ȋL$�D3T$�D3T$��E1�D�t$���ܼ���A��D	�D�T$��ω�D!�D!�	��������D։�����ܼ�D�T$�D3T$�	�A1�A1�D3t$��։�E1���D!�!�A��D3t$�	��D�T$�A�����D��D�T$�D΍�ܼ��Ɖ�E1�	�E1�D3T$�!�A��A����E���!�D�T$�D	�A��A��D�A�� ܼ�A��A	�E��A��A!�A!�D���E	�A��A��E�F��ܼ�E����E1�	�D3D$�D3D$�!�A��D�D$�A����D�T$�!���D	�E��D�A��D�D��>ܼ��|$�D��	�1�3|$�3|$�!��ǉ|$���D��A��!�	�D������|$��D��1ܼ��t$�D��D1�3t$�D1�D	��Ɖt$���D��A��!�D!�	�D�����t$��D��
ܼ��L$�D��D	�1�3L$�3L$����L$���D�ʋt$�D!�D!�A��	�D�����ʍ�ܼ�D�D$�D	ʉ�D��D1�3D$�D!�D!�3D$�	ʉ������B�A��3\$���ܼ���3\$�3\$�D	���D3|$�D3|$��щ���D3|$�D!�D!�A��	ʉ�E����B���ܼ���	�D!�A�҉���!�D	�A��A��D�A��ܼ�D�L$���D3L$�E1�	�A1�!�A��D�L$�A�щ�D�\$�!�D	�A��A��E���D�E��ܼ�D�D$���D3D$�D3D$�	�A1�!�A��D�D$�A�Љ�D�T$�!���D	�E��D�A��D�D��ܼ��|$�3|$���3|$�1�D1�D1�A���ǉ|$�D������|$������bʋT$�3T$�3T$�3T$����T$���D1�D1�����|$�A���D����bʋL$�3L$�D��3L$�D1�D1�1������L$�D���|$���D�T$�D3T$�ʍ/A1�D3T$�����b�D��A��1��D�T$�D1����D��A��D�T$�D�D����bʋL$���D1�D1�1�1�3L$����L$�D����ʋL$�D���D3T$�D�L$�D����b�D��E1�D3T$�1�D��A��E1�D1���D3L$�D3L$�A���D��A���D�T$��t$�D����bʉ�D1�D��D1����C�A��D�D$�����b�D��D3D$�D3D$�D1�D3D$���A��D1����A�8A���|$�D����b�3|$�D��3|$�3|$�D����D1���1�1�3t$���D1��B�D1�3D$�D����b�D����1�1�D����D1����B�.A��D����bʋL$���D1�E��1�3L$�D1�A��D1�D�A����A�E����b�D��D1�E��D1�A��D��3\$�A������bʋT$�D3|$�A��1�D��A��1�D1���D1�A��A�D�E��A����b�D�T$�E1�A1���E1�A��A1�A��A��E�E�G��3��b�D�t$�D3t$�E1�E��E��A1�A1�A��A��A1�E�E���G��5��b�D�t$�D3t$�E1�E��D1�A��A��A1���E1�A�A��E�G����b�D�d$�D3d$�D1�E��A1���A��D1�A��D1�D�A��D�A���bʍ�=��b�D��D1�A��A��D1�D�D�t$�D3t$�D1�L�D1���H�D���A��Dl$�D1�A��1�A��D�D�L$�D3L$���D1�L�1�D��DD$���1�|$�H�1���\$�A�D��D\$����IԋT$�3T$�1�A1�H�D$�A��M�D�XE�XD�(�xD�@H��[]A\A]A^A_�H�#Eg�����GX    H�H��ܺ�vT2H�G�����H�G�AVAUATI��UH��S�GXH����@uH�w�����CH���CX    �?H����   ��t4M��tHcCX��?�PH��I�̉SX�U��T��1�1�H������M��tgM��N�t% L��L)�I��?vH��I��@�����CX    �C��L��H��H��Hk��H��H�1�I�I9�tHcCX��?�H�KX�L H�L��[]A\A]A^�AUATI��USH��1�RH��1������CHcSX������Ѓ� D�,�    ����	ōB�CX�D���7HcCX��7?�P�SX�D ��HcCX��?�P�SX�D ��1�H��1�����H�S�   1�H���f��f�CP  A�H��f�kRH�kD�kTH�������ȉC�CȉC�CȉC �CȉC$�CCȉC(A$�C(A�D$X[]A\A]�H��κ   �t$H�t$����H���I��H���H��1��L��H��H�������SH����ZB 蹵����t0�K+$ ��%Hc¹2   H����Hi��   �,+$ H�f H���[��P�   ���B �I  H�?�' ZËD$�7�W�G    �GL�GL�OH�O �AWAVAUATUH��SH��H�GD�gD�/D�0H�G H� D��D�8D�@D�wE��y%A��u
�����A9�|A��u
�����A9�|D����D��A��A)́}�   ���B 1�D�D$�L$�ܯ��D�D$�L$�ERE��D��H���' P��X����  Y^���  tzD�m A�̅�uCH�E D��uD)�H��m  �2�ع
   E)��u�D��A������H�E Hc�H���C  ��tA���u�E��y!�uH��' H��A�}�[]A\A]A^A_�  H��[]A\A]A^A_�H�G�8 t�����H�D$�7�WH�G   L�GL�OH�O H�G0�U��SH��R��tH�G�8 tH�W0�w�?�  X��H��[]롉7�W�G����L�GL�OH�O �H�G�8 ��   H�WHcG���u9���   ����   AUATUSH��H�����taH�W D�'�oH���PD�(D�@A)��P)Ձ��   ���B 1�D�D$�1���D�D$PH���' D��E��U��X���D���  ZYH�C�s�;HcH�C H����  H�C� �CH��[]A\A]�É7�W�G    L�GL�OH�O �H�G�8 ��   H�G�O9u����   AWAVAUATUSH��APH�G �oD�'�PD�xfD�(fD�p)Ձ��   ���B 1��e���H�C�8 tH�S �s�;�/  �'D��RH��' A��UD)���X���E��A���(  Y^H�C� �CX[]A\A]A^A_��SH��   �1F  H�[�AVAUATU1�SH��H�����B �	   1�L�$�    H�|$�0��I��$�$f H�|$�Ӊ��B �	   H�|$1�H����/��I��$�$f H�|$��H��
u���$f �%�B 1��Ӊ�.�B �	   1�H�|$�/��H�4�@$f H��H�|$��H��uо�"f �7�B 1���I��M�>�B �	   H�|$I��1��a/��I��$`"f H�|$��H��$f H��I��$h"f H��u��sY$ �G�B 1�1�	   H�|$A��"f �/����"f H�|$�Ӿ0%f �N�B ��M��E1�E���T�B �	   H�|$1�A����.��L��H�|$I����A��uΉ�^�B �	   1�H�|$�.��I�t$H�|$�Ӊ�g�B �	   H�|$1��.��I�t$ H�|$�Ӊ�p�B �	   H�|$1��e.��I�t$(H�|$�Ӊ�z�B �	   H�|$1��A.��I�t$0H�|$�Ӊ麃�B �	   H�|$1����.��I�t$8H�|$I��@�Ӄ������ $f ���B �Ӿ($f ���B ��H��[]A\A]A^�SH���*D  H�    [Ã=�F$  tgRH�=:�' �G  H�^F$ 1�1��E  �=�X$  tH��C$ 1���   �)  �  H���' 1�1�PE1�A�    �@  h�   �   H���Ë��u.�G��f1ҁ�  ma��  = ema��  �F$    �u  X$ �i  USH��H���=�a$ u�s���e �������8  �  �w���e �������tVH��E$ ���   �у������   u)H�H��t
ǂ�   d   �@,d   Hǀ�   ��B �	  Hǀ�   ��B ��  �s� �e 莮����tWH�KE$ �  @1�H��H�H0Ǆ�      H��H��$u�H���   Hǀ�   ��B H���   H���   H���   �  �s�`�e �%�����tmH��D$ �  @1�H��H�H0Ǆ�      H��H��$u�H���   Hǀ�   ��B H���   H���   H���   H�      H�PPH�PXH�P`�  �s� �e 覭������   H�_D$ H�t$� �e Hǀ�   ��B �����D$�T$�=�}" t	�=�}" w��0k�
���S�|��)��1�����P~H� D$ Hǀ�   �B �   �|о   �   �u���# ����t�s�@�e �������u�U�s���e ������t*H��C$ ���   �у������   uHǀ�   �B ��&�# ����t�Hǀ�   .�B 1�Hk�H�sH��@�e 荬����tBH�=JC$ H���x8 u	���
���H��t	�@8   ��G<    H�C$ Hǀ�   C�B H��H��u��s���e �0�����tH��B$ Hǀ�   T�B �   �s���e ������t%H��B$ ǀ�      �@8   Hǀ�   ��B �Z�s� �e �Ы����tH���B �4   � f Hc�S$ Hi�H  H���;f �H8D�HD�@1�����H�WB$ Hǀ�    f �=�T$  ��   �S���H�t$���e ������{" �t$�T$��u��0k�
�Tо   ���0��0�=�{" 	t���W�   ��~N��u�����u�����u
��1��	���u
��"��(H��A$ �=I]$ Hǀ�   ��B ����H��1�[]�1��H��A$ �d   ���z,dNJ,9�# t)Ⱦe   �
�# ���������8$ ��8$ �R��8$ ��	��   H�5A$ �z, u#��8$ 	   �9$ )   �9$    �B  ��\���    tS1�1ɋ��   9�`f t��`f �   H��H��$u܅�t'�H8$    ��8$ F   �,�������8$ �M  �=$8$ ��   H��@$ ���    ��   H���   H����   H�:H9���   ��7$    �R,+c�# ��~�<8$ #   �������*8$ �P  �P�w�H��*���H�!@$ H��z89�s)�=   ���A���)ǁ�   �A����7$ #   E���\��������w����P��E��D�7$ �=C7$ cH��?$ ���    tS�@,+��# ��~�7$    �7$ #   ����������6$    �a7$ #   ��������O7$ �   �=�6$ lH�N?$ ���    tR��# ���u�Ԡ# F   �E�ȉʠ# u;��6$    ������6$    ���#    ����6$ �   ���# �����=b6$ 6H��>$ ���   u�x8 t �@6$    ��6$ (   ��6$    �:�=�6$  u1�����   �}6$    �6$     �ƋS6$ ����\6$ �Z6$ X�RH�`>$ � �e �A|H��Hk����_d ��tH����   � ;$ 1�H�5�:$ ����|�P ����E����|�\ �<�@f t��@f H��H��u�������Q$ �6$     �5DO$ H�=�=$ �����=�=$  �Љ�=$ ��!�����=$ 1�����!�1҉�=$ 1��L�l9�t��)�H��H��u��5$ �p=$ X�P�k=$ ������H5$ ����H�d=$ �@,�c�# Z�H�R=$ S�P<���   ��t�Ѻ   ��)�9�Lڅ�t���   ����O����;���   ��t���   ����O؃�	��@D�   =�   ����t�   �=hv" 	u�C����   F�9�4$ t)��4$ i�   �=�<$ �   �9  Hc�H�<[�uE  [�U1�S��R�p<$ �2P$ ��t1Ʌ������K<$ �޿ "f ��1�����1�!ȉ,<$ ����H��`f �������H���f ��H��0�����H���   u׉޿�!f �@ f �����޿ f ������޿`!f ����H���H��0�#���H��`!f u�޿  f �����޿`f �����޿�f ������޿�f �����X�޿�!f []�c���P��;$     ������   Z�����1�������   Q��t1��=r�#  ���Q;$ 1�5Y;$ ���P;$ ������=D;$  tZ�X븿0�A ����P��RB ��6  �;$ Z�⿣�A �������HcsL$ �;$    ��:$     Hi�H  ��:$    ��:$     ��2$     ��2$ ����H���;f �ǡ# ����H��:$ 1���d<f H����\f H��$u�H���H�t2$ �v2$ �����H��:$ ATA�H%f ��$f U�,   A�@ f �   S�B|1�W� "f Hk�j���_d L����   ��   ����H�3:$ AXA�H%f ��$f �Z   ��!f �P|�5�9$ L�@,��6$ ��   �����A�H%f A�@%f H�L7$ ��   �h   �`!f �����AYAZ��H��L��A�<%f �H��I��0��H��`"f ��k�
H��9$ k�L����   H�Á¬   ��o����H��u�P��$f ��   ��   jA�8%f A��f ��!f ����A�H%f A�Lf ��"f ��   ��   �  f �T���Z��$f ��   �5�8$ A�H%f ��   H�9$ � f L�@0�����A�H%f A�@f �@$f ��   ��   �`f �����A�H%f A�Df �@$f ��   ��   ��f �����A�H%f A�Hf �@$f ��   ��   ��f ����A�H%f ��$f H��8$ ��   �   �`f �$   L���   �����A�H%f ��$f H�S8$ ��   �   ��f �$   L���   ����A�H%f ��$f H�8$ ��   �   ��f �$   L���   �X���A�H%f ��$f H��7$ ��   �   ��f �$   L���   �$���A�H%f ��$f H��7$ ��   �:  ��f �$   L���   �����A�H%f ��$f H��7$ ��   �:  ��f �$   L���   ����A�H%f ��$f H�O7$ ��   �:  � f �$   L���   ������$f �:  H�7$ A�H%f ��   �0f �$   L���   �T���Y^[]A\Ã=��#  u%P�=�6$ �   �L3  H���?  �r�#    Z��R�=g�#  u����������!����L�#     X�P�^���1Ҿ   � (  �M6  H� �' Z�P轗��Z����SHc�Hk�H{6$ H�; t!�{詘����t�{荘��H��H(H�    [�AUI��ATUSAP�D�^E�U���vD)�A��A��D1�D)�E��A)�D����A1�A)�D9�B�, AO���)Ń=�Q$ t1���  ���   I��H�Ӊ�D��D���ƫ��A�U89�s)��������  ` �4���B ��������¸�   )Ё���� ��5$ A�$��H�=Q$ u(��  ��  �O�ȃ���  )����������  ���  )�������1��; ��Z[]A\A]Ë,�# H�15$ 1�9�~H�: tH9zu��������H�����AUATI��USHc�H����4$ �D$�C���lv�޿��B 1�覘��H��H��H��@ce H�z t!�D$B$�D$���i  ��4$ 9�~�T$M��t]Hc�E$ Hi�H  H���;f L9�tCH�T$L��H�L$�&���Hc�E$ Hi�H  H���;f H�rI9t$u�D$�   ��u��   �D$�   L��E1�������"�# H�'4$ A9�}$H�8 tM��tL;`u
D�������	A��H���׋�# A9�uAH��H�5�3$ 1�H��H��@ce A��9�~Hk�D�AH��H�<>D9G|��9�tlD���(���Ic�H��3$ H��Hk�H��@ce H�H�L�`�S(�ҍB�   H{, �C(yH���Ӕ���C,�L$�T$D��H��H-V3$ �?����EH��[]A\A]�H�=+3$  t�=*3$  uP袕���3$    Z��H�=3$  t�=3$  tP茕����2$     Z��AVAUATI��US1�H���X���9ϙ# A����   Hk�H-�2$ L�u M��t{�}������th��2$ I�~ �D$�   �D$tA�V$T$��~A9�}�D$H�uH��t7L9�t2L��H�L$H�T$����D���t�}�T$�t$�����������H���Z���H��[]A\A]A^�S����v��1����B �ߕ����[�x���S����v��1����B �������1$ [�U���@ce S��m   R�*����������������k=��# 1Ҿ   �i1  ���# 1�H��1$ 9�~Hk�H��H�0    ����1$     1�ǀ�ce ����H��@ǀlce ����H=   u�X�   [���A ]�F����.���H�=<1$  tOR�=:1$  t�Ó��� ���H�1$ H�x�Г��H�1$ �x�*.  H� 1$ H��0$     H�@    X��U��SH����u�KC# �����    F��G���Bv��1���B 1�舔���Hc�H��H���~e H9�0$ tj�O����{ u&H��'�B �	   1�H�|$�"���H�|$�!,  �C�{�   ��,  �{H�C�+,  H�{��������H�CH�������H�.0$ H��[]�S1�H��09�# ~Hk�H0$ H�8 t������H���ۋ�K$ �=zi" ��/$     �x t-H�|$�@�B �	   �=tC$ ��	�ύ<�����H��|�H��0�   [����1������   ���  v��    ��1ҿ   ��=   G��H�42$ H9�/$ u:AUA��ATA�ԉ�U����S����i P�R���YB�T-�B�t#���i []A\A]�7����AWE��AVLc�AUE��ATLc�U��SH��H�T$�\$PE��x9C�&=@  .��x*B�=�   E��xC�=@  ��xA�=�   ~���C 1�萒��D���D��D���6���i�@  Mc�i�@  Hc�Hc�I�L�.$ L�HT$E��~L��H��L��H��@  �I��@  A����H��[]A\A]A^A_�H�=q.$ �ATUH��S�B)��B��)�H�T.$ Lc�H��u�M D�EE��y�-��H��D���Ѕ�u��   A�=@  ��xB�=�   ~P�E��D��D�M���C P1�袑��ZY��i�@  �M�U D���>����} 1�Hc�L�H�-$ L�9�~KHcD�H�����t6Hi�@  D�H1�L�L9�tLi�@  D�\0H��F����PH�D��H���[]A\�ATUH��S�B)��B��)�H�R-$ Lc�H��uE��y�2��H��D���Ѕ�u��   �E D�=@  ��x�E�=�   ~��C 1�贐�����M�U i�@  D���R���L�E 1�Hc�L�J�|� H�,$ L�3A9�~NHcGH�����t6Hi�@  D�P1�L�L9�tLi�@  D�dH��F�$���PH�D��H��H���[]A\�����ATUH��S�B)��B��)�Lc�x�D�=@  ��x�B�=�   ~��C 1��ޏ��i�@  D�E 1�Hc�L�H,$ L�3A9�~dHcT�H��<�tPHi�@  �zL�RL��σ��t,�E�H@  I����D�L��+$ Hc�A����������BH�T�H���[]A\�ATUH��S�B)��B��)�H��+$ Lc�H��ui�@  D�E 1�Hc�L�Hm+$ ���H��D���Ѕ�u��nH��L�3A9�~bHcL�H��<�t�Hi�@  D�QH�yL�A��A���t,�D�H��H@  ��D�L��*$ Hc�A����������AH�L�[]A\�ATUH��S�B)��B��)�Lc�x�D�=@  ��x�B�=�   ~�,�C 1��K���i�@  D�E 1�Hc�L�H�*$ L�3A9�~dHcT�H��<�tPHi�@  �zL�RL��σ��t,�E�H@  I����D�L�,*$ Hc�A����������BH�T�H���[]A\�AWAVAUATI��USQ�B)��B��)�Hc�x��=@  ��x�B�=�   ~�A�C 1��u���i�@  L��)$ E�$1�Hc�À  Hc�H�H�DL�I�I�L�A9�~lIcL�L��<�tXHi�@  D�q1�1�M�,H�I9�t1D�8L�=L)$ A��Mc�G�D�8D�D)H��E�D= H��@  ���AH�L�H���X[]A\A]A^A_�P�   �Y�C ��%  H��($ Z�P�   �a�C ��%  H��($ Z�AVLc�AUA��ATM��UHc�S��E��xA�.=@  ��x
�=�   ~�h�C 1��P�����i�@  D���D�������Hc�L�H�($ A��A���tH��L��H��H��@  �I����[]A\A]A^�i�@  Hc�Hc�H�H�=�*$ H�1�9�}1�9�~	D�H����H��@  �����i�@  Hc�1�Hc�H�H5�*$ 9�~�H�����i�@  Hc�1�Hc�H�H5*$ 9�~Hi�@  H���>���SA��D��A��A�������C�t�D������D��D��D������A�|�D��[�H����>  H�=�'$ ���H�='$ �H�*$ H�p'$ �AWA��AVA��AUD��I���   ATA��1�UH��SC��6�  H��L�D$��&  �   L�D$H��H� 
A�D$�f�CH�SA�G�f�C
H��1�H�SFfD�cfD�{�H�׹:   �CAfD�cBH���   f�CD �1�A9�~+A�L �΃��@���t�
H�����A�L H���J�H�����1�A� �LH��H=   u�H��  H��H��H)��$���H��H��[]A\A]A^A_�E%  UH��S1�H��H��1�A�x�C ��H��   軺��H���e�����t�Ã�duӿ|�C 1��ŉ���   ��RB ��"  H�5�($ H���   I���@  ����H��[]�AW�w   �w   AVAUATUS���w   H����.  �U   �U   �U   �D$�.  1�1���   A���.  1�1�1�A���.  1Ҿ�   ��   A���.  ��   ��   ��   A���i.  �=�'$  �  ���# �q� �\I� TR� �Z�f/���   D�D$�	   �x   �ž   ��   �����	   E���x   �   ��   ������# 9�)��*��^�# �,��k�(A�w   �   ��   �ؙ��D��v   ��w��DN��������'D�¾   ��   �%�(   �   ��   �V���D��   ��   A�P��@���H��D��   [�   ]��   A\A]A^A_�@���H��[]A\A]A^A_�SH��   ��   H�[�AWAVAUATU1�SH��H��(�=_]" uJ9-�%$ ~/����C �	   1�H�|$��
��H�r$$ H�|$H�4�H�����ɾ�&f ���C 1����  H��%$ A����C �	   H�|$�1��}
��H�&$$ H�|$H�4�H����H��	uþp'f ���C �Ӿx'f ���C �Ӿ`'f ���C ��H��%$ �8�1�H��%$ A��l$Hc 9,�@�C �`���Lk�HL� �C E1�M��M�j E��E9f~OH�L%$ ���u�|$t%H�|$E�����C 1��	   ��	��L��H�|$���J�倏e I�E I��I���H���l������C �	   1�H�|$�	��H�4� 'f H��H�|$��H��
uоX'f ��C �Ӿ�&f ��C �Ӿ�&f ��C �Ӿ�&f �#�C �Ӿ�&f �*�C �ӿ1�C ��&f �ӿ9�C �#  ��x�=o4$  t�=�5$  u��&f �9�C �
��&f �?�C ��1��&f �F�C �ӾP'f �M�C �Ӿ�&f �U�C �Ӿ�&f �\�C �Ӿ�&f �d�C �Ӿ�&f �j�C �Ӿ�&f �r�C �Ӿ�&f �z�C �Ӊ麁�C �	   1�L�$�    H�|$�j��I��$`&f H�|$�ӍM���C �	   H�|$1�H���?��I��$@&f H�|$��H��u���Z" ��u�	   �TB H�|$�R����)H�b#$ �
��u��t׺��C �	   H�|$1�����H�|$�(&f ��H��([]A\A]A^A_�SH���  H�    [�H�T!$ 1�1��C���1��USH��8H��"$ �= Z" Hc@u9�"$ ~pH�'!$ �@  �   ��H���)Ɖ�   ���H�ʉ������H��"$ �   H��!$ HcPH�� $ H���P������p�)Éؙ��H�ʉ��}"H�|$���C �
   �H�T$�   1�����H��8[]�U�   S�@  PH�7!$ ���)Ɖ�   ���H�ʉ��T���H�"$ �   HcPH�M $ H���Q������p�)Éؙ��H��Y[]������H��!$ Hc�H��Hc H��H�H��<�`�C ��d�C D�BA��E)�D�E�A��?  &E��x!D�BA��E)�D�BE�A���   E��ySH�VH��t;�rA��A)��2DƁ�?  #E��x�rA��A)��rDƁ��   E��y�q���C 1��������R����=X" ��   H�� $ �8��   ATU1�SH�� $ Hc 9,�@�C ~gHk�HH� �C ��C@������u�� $ D�`荳����{���u�� $ �CD�d�o�����{D�S8���u�o $ ���C8H���[]A\�Ã=|W" ��   H�[ $ �8��   ATE1�USH�D $ D��HcD9$�@�C ��   Ik�HH� �C � $ 9S8u{���t!��t��t>�i�C@���C@;C|V�C@    �M�C@���C@;Cu@�C@����S��謲����{��*�=�$  u��t�C9Au�C@�H�K@;Ku�C@S�S8I���K���[]A\�Ã=�V" tMH��$ �8AS1�H�q$ Hc9�@�C ~)Hk�HH� �C HcP@��xH�T� �p�x����H����[��AWA��AVA��AUATA��U��SH��H�9$ D�(��y��t+��1�
   �������u�D��1�����D1�)��  u	�l1ҽ   ��E���˃��t7�й
   E)�D���D��D�L$��Hc҉D$H�� 'f ������T$D�L$��A��D��)�E��y��H��$ D��������H����[]A\A]A^A_Å�x*ATA��H��$ U��S������D���߃��[]A\�����Å���   AVAUA��ATA��U��S��  ]�   A�<   D��   ��D����k�<�A������H�X$ �)ЉŃ�<t
D�������t2H��D�������D�������u��H�z$ []A\�A]A^)������[]A\A]A^����$ ������$     �l$ 
   �Q�����_$ uZ�_��X��_$    �]$     �7$ �   �,���Q������&$ �ȉ$ t	�=1$  tZ놃��������N$ X�USQ������k����=T" uH��$ �xu�~H��$ �8~Z[]�����X��u�X��1�9���`'f ���������H��$ �x t�`'f �   �����=�$  tH��$ �p'f �x�����=�S" u��s���X[]���$    �J���Hc�1�1�Hk�(H8$ �<��9f  t9�tD�H��H��u�+D���$     1��$     �@$    ��$ #   ���9f  t2H��    1҃��9f  tǄ�%f     H��H��u�ǀ�%f     H��H��u�����S�7����=�$  ��   �=�$ t|��$     L�w$ E1�B�<��9f  D��t;Ik�(L��1�H��Lʃ��9f  t�t���%f H��H��u������B���%f I��I��u��R   1������T$    �N$ ����   ��$ u�   1��y���L��$ E1�E1�B�<��9f  D����   Ik�(L��1�H��H�%f Lփ��9f  t:D��\A9�t.A�K��yA�K���c~� c   ����|��� ����A�   H��H��H��u�������c~B���%f c   ����|
B���%f �B���%f ����I��I���G���E��ua�R   1������S$ �M��u*�=$  t?1��   �����=Q" u[�R���[�����t��$ u�x$ #   ���$ [�AWAVAUATU�   S1�R�������������   �  H�@$ f���f��f��H�ʾ-   �)������d   �
   H�#$ �����2   �   H�$ ����Dk�!Dk�(A��DA��R�<��9f  ��   H��`&f D���#   A�*   f���f��f��H�ʘ)��=���H��`&f D��D��f���f��f��H�ʘ)�����9�$ uTH��`&f D���#   f� ��f��f��H�M$ �)������H��`&f D��D��f� ��f��f��H�,$ �)�����H��H���'���H��$ 1�D�(E�uRDk�!A��N�<��9f  tRI��1�I�����9f  tk�
A��/�%f �   D��D������H��H��uҋ��%f A��  �   D�������H��H��u�X[]A\A]A^A_�RE1���$     ��$     ��$    �e$ #   B�<��9f  tDB���%f     D��B���'f     B���'f     B���'f     �$���8$ �2$ I��I��u�1��= $  ���$ X�7���V������=L$  ��   �=�$ 
��   H�$ L�$ E1��$     D��$ L�HB�<��9f  tJAkd�A�zB���'f AkAd�A�zB���'f AkAd�A�zB���'f E��tD���d���B���%f I��I��(I��u��R   1������O$ 
   �I$ ��uk�i$ u�   1������L�\$ L�]$ 1�1����9f  t/���'f �pHk�
���'f AkDd�A�x9�|���'f ��   H��H��u��n��u{��$ u�   1�����L��$ L��$ 1�1����9f  t/���'f �pHk�
���'f AkDd�A�x9�|���'f ��   H��H��u��R   ���o  �  ����   �u$ u�   1�� ���L�h$ L�i$ 1�1����9f  t/���'f �pHk�
���'f AkDd�A�x9�|���'f ��   H��H��u�����   1��R   �����=�$ ������$ ��   ��uy��$ u�   1��e���E1�E1�B�<��9f  t1B���%f D��D�HF���%f �]���A9�|
B���%f �A�   I��I��u�E��ua�9   1��	����>$ �M��
u*�=|$  t?1��   ������=kK" uY����Z������t��$ u��$ #   ����$ X�AWAVAUATUS�   RH��$ �(������u���� ���H��$ �2   H��$ f� ��f��f���=�$ ҃� ��|`�H��)�����H�d$ �2   H��$ f� ��f��f���=e$ ҃� ����   �H��)������H�$$ �2   H�`$ f� ��f��f���=%$ ҃� ����   �H��)������=$  t3H��$ H�$ �2   f� ��f��f��H�ʘ��   �)��G���H��$ 1�A�   D�hA��2�<��9f  ��   H��$ D��f� ��f��fA���=�$ ҃� �D�d H��`&f D���)������9�$ uH��`&f D��H�1$ D��� )�����E�u
���'f A�|$@)�D����������'f A��$�   D��)���������'f A��$�   D��)�������=�$  t���%f A��$   ���D�������A��!H��H������X[]A\A]A^A_���$     ��$     ��$    ��$ ������$ ������$ �����Z$ �����T$ �����B$ #   ����V�����=�$  ��   �=7$ 
��   Hcv$ 1�H�5a$ �g$     Hk�(HD$ kAd��~�$ kAd��~� $ kAd��~��$ �A�#   �����$ �F �R   �����$ ������$ 
   ��$ ��uQ��$ ��$ u�   1��S���Hc�$ H�=�$ Hk�(H�$ k@d��9�$ ��  �w$ �T��uf�Y$ �r$ u�   1������Hcy$ H�=f$ Hk�(HS$ k@d��9$ �@  �$ �R   1�������$ �#  ��uQ��$ �$ u�   1�����Hc$ H��$ Hk�(H�$ k@d��y9�$ ��   ��$ 듃�u{��$ u�   1��C����h$ �#   �pHc�$ Hk�(H�$ �@���9Ɖ�M��7$ �55$ �pH�w$ �5!$ �@ ���9�|`;$ �$ R������
u*�=X$  t?1��   ������=GF" uY����Z������t��$ u��$ #   ����$ X�U�   SVH�$ �@�@�����������k2�\2�I���������2   �2   H��$ �������$ �2   �  �D���H��$ ��2   ������`$ ��  ����H�}$ �޿2   �����+$ �޿  �������   �   H�&$ ������$ ��   ��   �����H�-$ �8.H��$ ��   ��   �R�����$ ��   Y�0  []�����X[]Ë $ 1�1ɸ�;f @�A�   �<��9f  tXD�HA��t���    ǀ�      D�AD��
ǀ�       A��t���    ǀ�      D�AD��
ǀ�       H��HH  H��u���t�s$ �AQ�J$ ���B$ ��u�=[D" �   �C   t�   ������6����.$ ��t��t/��u1Z�����=<$  tAX�W����=�$  t_����^�]���Y����X�R�=�C" u1Ҿ   �   �n$     �1Ҿ   �H   ��	  �hB H��
$ �=����   ���C �"  �   ���B H�*$ �  H�$ Xÿ�B ������j$ ��t��t*��u+������=y$  t�����=;$  t�����*����"���ËG$� H�=$ �!$     �$ H�G(��$     ��$     H��$ u�G   � u�G   � u�G   �=�B" t���~����V����������=�$  tY�y����=�$  tZ����X����AWAVAUATU1�SH��   H�|$H�|$$螹���p$     9-z$ ��   ��	   H�|$Hk�(Hu�' H������H�|$$H�t$����L�kD�5+$ 1�H�=*$ ��A9�~H��L;l��u��)E�~Mc�I��L���d���D�=�
$ D��H��
$ N�l �H�|$$�������sH�|$$������sH�|$$�����K���H�|$H�t$$�޹��H�Ĉ   []A\A]A^A_�SH�����C �p��H��H�:v# [��H��`H��`AT�   ���C US�=p����1���tKHc�H����9-q&$ t5H�p&$ H��H�<�?-t!�
���WB I��H��1�����L���B   ���   []A\�ATI��U1�S�  A�<,@��t�c�����H����1�1�H��u߉�[]A\�AWAVAUATUSH��H��(�"���I��H��uH�޿��C 1��=����  H���1�H�߾/PB �-�	$ H��H�|��U�����t71Ҿ   �   ���  H��I���     A�EI�t$A�D$�ٖ���   1�H�T$L��   �����   ���C H�|$�������t'�   ���C H�|$�������tH�޿��C 1��6j���\$1Ҿ   �����  �t$Hc�L��H��I���L���l$Hc��(   D�5�$ ����H��H��u���C 1���i��H��E1�D9=�$ H�=��' vzA9�suIk�(�
   H�4H���H�zH��tH�rH�D$H�$�	  H�D$H�$H�i�' H�D H��t"H)�H���������H��H��H�Hk�(H�H�B I��H��(�v����l���IcƉ-$ M�|$Hk�(H��' H�A9�s7A�G�L�kL��H�ߺ   H��(A��I���C�A�G�H�C�    �C��f�����L���'  H�=�$ H��t�  H��$     H��(L��[]A\A]A^A_Ë�$ �ATI��UH�-z$ S�k$ H��tC�I���1���Hc�H�\� H��t]�   L��H��������uH+M�' H��i������9H�[ ����Hc�Hk�(H-+�' ��xH��   L��H��(�c�����t���������[]A\�UH��SQ�_����Å�yH����C 1�� h����Z[]�S��9�$ w�޿�C 1���g��Hk�(H��' �C[�9=�$ ATI��U��Sw��1��)�C �g����Hk�(H��' �E  HcK�sL��H�{������S9�~�Ɖ�D�C 1��vg��[1�]A\�  AUA��ATA��USQ;=!$ r��1��n�C �Hg��Ic�Hk�(H�' H�CH�hH��t	HcCH��IH�kH��t��  ���C D��H���0  �)D������H�SD�����  D��H�CH������H�kZH��[]A\A]�H���t$�����t$H�����I���SHc�;s$ r�޿��C 1��f��Hk�(Hp�' H�CH�x uH�{��  ���C [�   �  [�P�C���Z���AUATUSRH�=!$ H��t�  �=	$ ��tc��1Ҿ   1��  ��$ I��H��$ 1�H��L���D�-�$ A9�v+Hk�(Hڕ' H��H������1�A��I��H�H�S H���X[]A\A]�AUATA��US1�H����`�C D9�tSH��h�C �������xC���!��D��H�D$�!���   ��I�����A���C L�L$L��H��L�¿��C 1��de��H��H��@u�H��[]A\A]�H�G8H�H�G(H�G H�G0H�GH�GPH�GX��G   ��8�GH   �G8�H��H�|$�Bg���T$H�H8H��' H�H(���8H�H H�H0H�HH�@�@   H�HPH�HX�@H   �P8H���UH�o�SH��R��J t���C 1��d���{�tH�C�H��tH�     H�C��C�   H�C�    �x�C�    u$�S�H�S�H�PH�B H�@�' H9j0u	H�B0�H��H�P�zu!�
H�JH�HH�A H��' H9Q0uH�A0X[]�AW��I��AV���AUA��ATD�g(USQH���' H�h0H�E �xHD�L�u H��L9�uD����C 1���c���E��t%��	H�mH���H�[ H�}(�����H�[H�k�H�m�{u��D9�|�D)��@~.Ic�H؉H�S�@   H�@    H�X H�PH�B H�CD�#M��uA��~���C 1��Ac��L�{H�C(D�kM��tI�H�KH��' H�J0�CJ Z[]A\A]A^A_�H��' ATU��S��H�x H�ڒ' H��H9�t(�GL�g9�������t9�	H��(����L����[]A\�H���' ATA��U���%�C S�0H��1������D���B�C 1������H�k�' H�X D�CE9�A9�|H�K�H�޿W�C 1�����H�=�' H�SH��H9�tIHcH�H9�t
���C ����H�CH9X t
���C �o����{uH�C�xu
���C �U���H�[�[]A\�U�%�C H��SRH�Б' �H��1��|���H���' H�X D�KL�CH�ھW�C �H��1��U���H���' H�SH��H9�tUHcH�H9�tH���C �i���H�CH9X tH��7�C �R����{uH�C�xuH��h�C �5���H�[�{���X[]�H�)�' SH�X H��' H�SH��H9�tOHcH�H9�t���C 1��a��H�CH9X t���C 1���`���{uH�C�xu���C 1���`��H�[�[�AUA��ATI��U��SH��AP��J t��L��$�C 1��`����~H�{� uD��L��P�C 1��`���k�X[]A\A]�UH��SH��R��J t���C 1��b`��H�k�H�] X[]�H�8�' 1�H�Q H��H9�t�r��t��~H�R���H��' � �AT��I��UH��1�SH��H�����H�KL��[H��   ]A\����SH��H�����H��[����U�P�B SQ�,���H��1�H��t51Ҿ   �    ����H��H� ��e H��H�@    �]���H�k�CH��Z[]�H��(H�t$H�|$��  ����   �T$�L$�Ѕ�t���u�   ����uM���5�# ��t;�=�#  �D$    �T$~��xHc�����C �1��D$��t�H�|$�#���끺�   �D$   �T$�D$    ��t
H�|$�����H��(�Ã=fi#  �    IZi# E1�H�L� D9�~?F�I��J��@(f �A�I����������	�B��@(f ����	�f�L���E1�A�   D9��SB�D��+r$ H��@(f D�HD�@A���S$ E��A��D��+O$ A���B$ A��D��@(f ��D��+6$ A���)$ A	�A����D	�E1�D9�h# ~2E1��� $ J���D9�vB��    ����B�I����A��H����I��D9��G���[ù�  ��  �`�C H��  �  RA�    A��  ��  H�{ $ H�| $ �  ��� $     H��H�j $ H�      H�a $ H�      H�` $ 1��L $    �R $    �m����C $ ���C D� $ D�4 $ � $ Q�5 $ � $ P� $ P���# P1��+���H�� �@  1��!�C ��   �����   �S�C �Ga����~"H��$ H�H�|�������\�C �$g# ���0���# �@  1ҿ��C ��1ҹ�   �Ƌm�# ��9�G��5�f# 1�����1Ҿ   � �  �*����=>�# �=;�# H� �# �:�# ����������'    H���# X�.���PH�=��# �6���H�=��# Z������_����AWAVAUATUSQ���# L�5��# H�-��# iRf# @  M�� �  )��# ��A����A��D)���M9�tHE1�D9="f# ~3L�@  L��A��H����������# ����e# i�@  �H���I��@  볋Z�# H�5+�# 1�H�=r�# ���0�# ��e# i��   �Z[]A\A]A^A_��  H�5��# ��>  ��Hc��# 1�H��H��B Hc�H������C(f  �w�@�40@�4�B(f �w�@�40@�4�A(f �w�@�40@�4�@(f ��   u��ATA��UE���S�����C �������1ɾ���1�D�+9�~�։ȅ�t
����   u�[]A\����  ������P� � ����H�u�# 1�Z�   S��   ����ztz��w��tqw��
t;�0�� t;��xt=�$��  t:w
��
  t7���  t4��  t3��������/�   �(��   �!��   ���   ���   ���   ���   �t�# ����	�[H��f��	 -f ���U�# �P���C ��,f H�2 2 ��H���# ������,f ��  � -f �   H��# H��1��Z�H��8H�|$�
  H��tAH�D$H��tH��tH��uۋt$ �   ��t$ 1��������H�=��# �h  1�����H���# H�5�# � � H���   ��  H�=��# �  H��8�1�Si�@B �'   �щ։��i[�S1Ҹ   �։�H�\$�H�L$��iiD$��  D$�[ËC�# 1�;?�# t!����f��  -f ���$�# �ԉ��   �SH��# H��tH��H�{,�����H��[��  [�UH��SH�}�L�E�H�M�   �    �    �    L���iH�E�[]�UH��SH�}�H�E H�E�H�E(H�E�H�E0H�E�   L�E�H�M�H�U�H�u�    L���i�[]�UH��H�}��u�H�U�H�E�H�P�H�U�H������tH�E��U�H�E��ڐ]�UH��H��0H�}�H�u�H�U�H�E��H��t(H�E�H�P�H�U�H������toH�E�H�U�H�H�E���H�E؃�H�E�H�E�H+E�H�E�H�E�H��H��H�M�H�E�H��H���  H�E�H�P�H�U�H������tH�E�H�U�H�H�E��ؐ��UH��H��0H�}�H�u�H�U�H�E��H��uH�E���H��tH�U�H�M�H�E�H��H�������   H�E؃�H�E�H�E�H+E�H�E�H�E��H��uH�E���H��t H�E�H��H��H�M�H�E�H��H����  �H�E�H��H��H�M�H�E�H��H���  H�}� t'H�U�H�E�H�4H�U�H�E�H�H�E�H��H���c�����UH��H�� H�}�(   �;���H�E�H�E��@    H�E��PH�E���E��H�E��P�E��H�E��P�E��H�E��P�E��H�E��PH�E�H�U�H�PH�E���UH��SH��H��H��H�M�H�]�H�U؋U؋E�9�|/�E؋M��U��9�} �U܋E�9�|�E܋M�U��9�}�   ��    []�UH���E��E��,��E��*E�f/E�v�E�����E�]�UH��H�� I��H��L��L��H��H�u�H�}��U�H�M��M��U��u�E�L�E��}�M��A�����  ���UH��H��@�}܉u؉UԉM�D��D�ɋE�ỦʈUȈEă}� y�E�E��E�    �}� y�E�E��E�    �E������E���	��E�	�   ��E�H�EH�@H�E��E�    �E�;E���   �U��E��H�E�@9�}u�U��E��H�E�@�E�U܋E��H�E�@9�|H�E�@+E���EԉE�}� ~,�E�HcЋM܋E�ȉ�H��    H�E�H��E���H��������E��l������UH��H�� �}��u��U�M�D�E�L�M��E����E�D���E�D���M��U�u��E��u�W������H�����UH��H��P�}̉uȉUĉM�L�E�L�M�H�E�H�H�UҋP�U��@f�EދE܉�HE��E��E��Eă��P��H����*��������E�E����E��E��E�    �E�   �E�    �E�;E���  �U�E��H�E��@9���  �E�    �E�;E��k  �U��E��H�E��@9��T  �E������E��E�Љ�H�E�H�� <uT�E������E��E�Ѓ���H�E�H�� <u,�E������E��E�Ѓ���H�E�H�� <��   �UȋE�Љ�H�E��@�E��ЋM̋E���E�ЉE��E������E��E�Љ�H�E�H�H�E�H�P�E�H����E������E��E�Ѓ���H�E�H�H�E�H�@�U�����H����E������E��E�Ѓ���H�E�H�H�E�H�@�U�����H������E������E�)E��E��E�E��E��F������UH��H��0�}�u�U�M�D�E�D�M؃}� y�E�E��E�    �}� y�E�E��E�    �E�    �E�;E��  �U�E��H�E�@9���   �*M��E����*��E����*��\��*U��^��Y��E����*��X��,����*M��E����*��E����*��\��*U��^��Y��E����*��X��,�D���*M��E����*��E����*��\��*U��^��Y��E����*��X��,����U�E��<�U��E��uQE��A���Ѻ   �������H���E���������UH��H�� I��H��L��L��H��H�u�H�}��U�M�L�E��M��U��u�E�D�E�}�H���u�E��A�����   H�����UH��H��0�}�u�U�M�D�E�D�M؃}� y�E�E��E�    �}� y�E�E��E�    �U�E��H�E�@9�~H�E�@+E���E�E��E�    �E�;E��  �U�E��H�E�@9���   �*M��E����*��E����*��\��*U��^��Y��E����*��X��,����*M��E����*��E����*��\��*U��^��Y��E����*��X��,�D���*M��E����*��E����*��\��*U��^��Y��E����*��X��,����U�E��4�U�E��uQE��A���   ������H���E���������UH��H��0H�}�H�u�H�U��E�    H�E��@9E���   H�E�P�E�)�9E���   �U�H�E��@�H�E�@9�~H�E�P�E�)��H�E��@�E��E���H�H�U�H�JH�U��R�U���Hc�H�4H�U�H�JH�U�RD�E܋}�D����U����Hc�H�H��H�������E��E������UH��H��@H�}�H�u�H�U�H��L��H��H�E�H�UȋU��E��H�E��@9�~H�E��P�E�)���EȉE��UċE��H�E��@9�~H�E��P�E�)���ẺE�U؋E��H�E�@9�~H�E�P�E�)���E��E��E�    �E�;E���   H�E�P�E�)�9E�}v�E���H�H�U�H�J�uċU��H�U��R����Hc�U���Hc�H�H�4H�U�H�JH�U�RD�E܋}�D����U����Hc�H�H��H��������E��k������UH��H�}�H�u�H�U�H�E�H�@H�E�H�E�H�@H�E��E�    H�EЋ@9E���   H�E؋P�E�)�9E���   �E�    H�EЋ@9E���   H�E؋P�E�)�9E���   H�EЋ@�E��E��H�H��    H�E�HЋ ��=�   vWH�EЋ@�E��E��H�H��    H�E�H��ŰE��H�E؋@�ЋE�E��H�H��    H�E�H����E��I����E������]�UH��SH�}�L�E�   �    �    �    �    L���iH�E�H�@tH�E�H�E�[]�UH��SH�}�H�u�H�U�L�E�   H�M�H�Uо    �    L���iH�E�H�@tH�E�H�E�[]�UH��SH�}�L�E�   �    �    �    �    L���i�[]�UH��SH�}��u�L�E�   �M�    �    �    L���i�[]�UH��SH��XH�}���   ��	  H��H�޸    �   H��H���H�H���  H�]�H�E�H���   H�E�H���   H�E�H��H�������H�E�H�E�H�U�H�PH�E�H�H H�E��|   H��H���s���H�E��@���E�H�E��@���E�H�E�H���   H�E��E� H�E�H�U�H�M�H���   H���   H�U�H�M�H���   H���   H�U�H���   H�E�H��X[]�UH��SH��H�}�H�E�H�@H������H�]�H��tH���  ��   H���	  �H��[]�UH��SH�}�H�E�L�@H�E�H�P �   �    �    �    L���i�[]�UH��H��H�}�H�E�H���   H�E�H���   H9�u-H�E�H���   H�E�H���   H�E�H�@�   H�������+H�E�H���   H�E�H���   H�E�H�@�   H����������UH��H�� H�}�H�E�H���   H�E��@&��H�E��@$��H�M苉�   I��A�ȉщ¾    �    �����E�    H�E�H����  9E�����t0H�E�U���H����  H�H�H�M�H���   H��H���҃E��H�E�H���   H��tH�E�H���   H�U�H�    H����H�E�H���������UH��H��0H�}�H�u��E�    H�E�H���G  9E�����t{H�E؋U���H���>  H�PH�@H�E�H�U�H�U�H�M�H�E�H��H���������t6H�E؋U���H���  H�H��H�H�M�H��H����H�E؋U����   �	�E��o������UH��H��H�}�H�u�H�E����   ��xLH�E����   ��H�E���H���!  H�H��H�H�M�H��H����H�E����   ��H�E���H����  �H�E�ǀ�   �����    ��UH��H��0H�}�H�u�H�E�H�U�H���   H�E؋��   ��x5H�E؋��   ��H�E؉�H���  H�H�� H�H�M�H��H�����   �E�    H�E�H����  9E�����tnH�E؋U���H����  H�PH�@H�E�H�U�H�U�H�M�H�E�H��H���_�����t)H�E؋U���H���  H�H��H�H�M�H��H�����	�E��|������UH��H��H�}�H�u�H�E�H�U�H��H���  ���UH��H�}�H�E�f�   H�E�f�@  H�E�f�@  H�E�f�@  �]�UH��H��H�}�H�E�H���   H�E�H�@    H�E�H�� H������H�E�ƀ�   �H�E�ƀ�   �H�E�ƀ�   �H�E�ƀ�   �H�E�ǀ�   ����H�E�Hǀ�       ���UH��H��H�}�H�E�H���2   ��ÐUH��H�}�H�E�H�     H�E�H�@    H�E��@    �]ÐUH��H��H�}�H�E��@��tH�E��    H���  ���ÐUH��H�}�H�E��@]ÐUH��H�}�u�H�E�@��tH�E�@9E�sH�E�H� H��uH�E�H� H�@�KH�E�H� H�E��E�    �E�;E�s)H�E�@9E�sH�E�H� H��tH�E�H� H�E��E���H�E�H�@]�UH��H��H�}��u�U�H�E���H���X�����UH��H�}�H�E�H�     H�E�H�@    �]�UH��SH��(H�}�H�uп   �  H��H�    H�C    H�C    H������H�]�H�E�H�     H�E�H�@    H�E�H�U�H�PH�E�H� H��uH�E�H�U�H��,H�E�H�@H��tH�E�H�@H�U�H�H�E�H�PH�E�H�PH�E�H�U�H�PH�E؋@�PH�E؉P�H��([]�UH��H��0H�}؉u�H�E؋@��tH�E؋@9E�r	H�E���   H�E�H� H�E��E�    �E�;E�s)H�E؋@9E�sH�E�H� H��tH�E�H� H�E��E���H�E�H�@H�E�H�E�H� H��t H�E�H�@H��tH�E�H� H�U�H�RH�PH�E�H�@H��tH�E�H� H��tH�E�H�@H�U�H�H��}� uH�E�H�H�E�H�H�E؋@�P�H�E؉PH�E؋@9E�����tH�E�H�PH�E�H�PH�E�H������H�E���f�     UH��H��H��H��fof H��H����H��]�UH��H��H��H���o� H��H����H��]�UH��H��H��~2fHn�f��f��fs�f��fs�f��fs�f��fH����H��]�UH��H��H��L��H��~ fHn�f��f��fs�f��f H����H��]�UH��H��H�}�H�}� uH�E�   H�E�H���������UH��H��H�}�H�}� uH�E�   H�E�H��������UH��H��H�}�H�E�H���b������UH��H��H�}�H�u�H�E�H����������UH��H��H�}�H�E�H���(������UH��H��H�}�H�u�H�E�H���	������fD  H��" H���t3UH��S�8Yd H��D  ��H��H�H���u�H��[]�f.�     �������                         Starting D_DoomMain AMMNUM%d Follow Mode ON Follow Mode OFF Grid ON Grid OFF Marked Spot %s %d All Marks Cleared fuck %d      p   `   @   �                             
               are you sure you want to
quit this great game? you want to quit?
then, thou hast lost an eighth! don't go now, there's a 
dimensional shambler waiting
at the dos prompt! get outta here and go back
to your boring programs. if i were your boss, i'd 
 deathmatch ya in a minute! look, bud. you leave now
and you forfeit your body count! just leave. when you come
back, i'll be waiting with a bat. you're lucky i don't smack
you for thinking about leaving. please don't leave, there's more
demons to toast! let's beat it -- this is turning
into a bloodbath! i wouldn't leave if i were you.
dos is much worse. you're trying to say you like dos
better than me, right? don't leave yet -- there's a
demon around that corner! ya know, next time you come in here
i'm gonna toast ya. go ahead and leave. see if i care. -iwad IWAD file '%s' not found! -iwad not specified, trying a few iwad names Trying IWAD file:%s
 unknown.wad Unknown game? Doom II plutonia.wad Final Doom: Plutonia Experiment tnt.wad Final Doom: TNT: Evilution doom.wad DOOM1.WAD Doom Shareware chex.wad Chex Quest hacx.wad Hacx freedm.wad FreeDM freedoom2.wad Freedoom: Phase 2 freedoom1.wad Freedoom: Phase 1 heretic.wad Heretic heretic1.wad Heretic Shareware hexen.wad Hexen strife1.wad Strife                         �OB           $OB     ,OB           9OB     YOB           aOB     |OB            I[B     �OB             �OB     �OB            �OB     �OB           �OB     �OB           �OB     �OB           �OB     �OB             PB     PB           PB     &PB            3PB     EPB           OPB     UPB           aPB     Disconnected from server in drone mode. Disconnected from server. TryRunTics: lowtic < gametic gametic>lowtic -testcontrols ENDOOM mouse_sensitivity sfx_volume music_volume show_messages screenblocks detaillevel snd_channels vanilla_savegame_limit vanilla_demo_limit show_endoom chatmacro%i PLAYPAL M_PAUSE  WARNING: You are playing using one of the Doom Classic
 IWAD files shipped with the Doom 3: BFG Edition. These are
 known to be incompatible with the regular IWAD files and
 may cause demos and network games to get out of sync. TITLEPIC demo1 CREDIT demo2 HELP2 demo3 demo4 titlepic INTERPIC MAP01 E1M1 E4M1 E3M1 -pack doom2 tnt plutonia Valid mission packs are: 	%s
 Unknown mission pack name: %s Unknown or invalid IWAD file. FREEDOOM FREEDM Unknown The Ultimate DOOM DOOM Registered DOOM Shareware DOOM 2: Hell on Earth DOOM 2: Plutonia Experiment DOOM 2: TNT - Evilution Emulating the behavior of the '%s' executable.
 Doom Generic 0.1 Z_Init: Init zone memory allocation daemon.  -nomonsters -respawn -fast -devparm -deathmatch -altdeath Development mode ON. -turbo turbo scale: %i%%
 V_Init: allocate screens. M_LoadDefaults: Load system defaults. doomgenericdoom.cfg default.cfg Game mode indeterminate.  No IWAD file was found.  Try
specifying one with the '-iwad' command line parameter.
 W_Init: Init WADfiles.  adding %s
 -gameversion 	%s (%s)
 Unknown game version '%s' dmenupic BFG Edition: Using workarounds as needed. -playdemo -timedemo %s.lmp Playing demo %s.
 
You cannot -file with the shareware version. Register! 
This is not the registered version. SS_START  WARNING: The loaded WAD file contains modified sprites or
 floor textures.  You may want to use the '-merge' command
 line option instead of '-file'. FF_END  WARNING: You are playing using one of the Freedoom IWAD
 files, which might not work in this port. See this page
 for more information on how to play using Freedoom:
   http://www.chocolate-doom.org/wiki/index.php/Freedoom I_Init: Setting up machine state. -skill -episode -timer -avg -warp -loadgame M_Init: Init miscellaneous info. R_Init: Init DOOM refresh daemon -  
P_Init: Init Playloop state. S_Init: Setting up sound. D_CheckNetGame: Checking network game status. HU_Init: Setting up heads up display. ST_Init: Init status bar. map01 -statdump External statistics registered. -record Supported game versions: Doom 1.666 Doom 1.7/1.7a 1.7 Doom 1.8 Doom 1.9 hacx Ultimate Doom ultimate Final Doom final Final Doom (alt) final2 chex                            �6@     7@     7@     47@     �6@     d7@     k7@             e2m1    e2m2    e2m3    e2m4    e2m5    e2m6    e2m7    e2m8    e2m9    e3m1    e3m3    e3m3    e3m4    e3m5    e3m6    e3m7    e3m8    e3m9    dphoof  bfgga0  heada1  cybra1  spida1d1        CTB            ITB            MTB                            [B     [B            [B     %[B            )[B     .[B            2[B     7[B            �OB     ;[B            @[B     N[B            W[B     b[B            h[B     y[B            �OB     �[B     	                               none heretic hexen strife                       }YB     CTB     ITB     MTB     �[B     ;[B     �]B     �]B     �]B                                                                    	      
                                                             	             	             	                                                                 	            	            	            <            "   Player 1 left the game -left -right -longtics -solo-net NOTE: Turning resolution is reduced; this is probably because there is a client recording a Vanilla demo. startskill %i  deathmatch: %i  startmap: %i  startepisode: %i
 player %i of %i (%i nodes)
 Austin Virtual Gaming: Levels will end after 20 minutes Levels will end after %d minute BOSSBACK PFUB2 PFUB1 END0 END%i VICTORY2 ENDPIC ZOMBIEMAN SHOTGUN GUY HEAVY WEAPON DUDE IMP LOST SOUL CACODEMON HELL KNIGHT BARON OF HELL ARACHNOTRON PAIN ELEMENTAL REVENANT MANCUBUS ARCH-VILE THE SPIDER MASTERMIND THE CYBERDEMON OUR HERO FLOOR4_8 Once you beat the big badasses and
clean out the moon base you're supposed
to win, aren't you? Aren't you? Where's
your fat reward and ticket home? What
the hell is this? It's not supposed to
end this way!

It stinks like rotten meat, but looks
like the lost Deimos base.  Looks like
you're stuck on The Shores of Hell.
The only way out is through.

To continue the DOOM experience, play
The Shores of Hell and its amazing
sequel, Inferno!
 SFLR6_1 You've done it! The hideous cyber-
demon lord that ruled the lost Deimos
moon base has been slain and you
are triumphant! But ... where are
you? You clamber to the edge of the
moon and look down to see the awful
truth.

Deimos floats above Hell itself!
You've never heard of anyone escaping
from Hell, but you'll make the bastards
sorry they ever heard of you! Quickly,
you rappel down to  the surface of
Hell.

Now, it's on to the final chapter of
DOOM! -- Inferno. MFLR8_4 The loathsome spiderdemon that
masterminded the invasion of the moon
bases and caused so much death has had
its ass kicked for all time.

A hidden doorway opens and you enter.
You've proven too tough for Hell to
contain, and now Hell at last plays
fair -- for you emerge from the door
to see the green fields of Earth!
Home at last.

You wonder what's been happening on
Earth while you were battling evil
unleashed. It's good that no Hell-
spawn could have come through that
door with you ... MFLR8_3 the spider mastermind must have sent forth
its legions of hellspawn before your
final confrontation with that terrible
beast from hell.  but you stepped forward
and brought forth eternal damnation and
suffering upon the horde as a true hero
would in the face of something so evil.

besides, someone was gonna pay for what
happened to daisy, your pet rabbit.

but now, you see spread before you more
potential pain and gibbitude as a nation
of demons run amok among our cities.

next stop, hell on earth! SLIME16 YOU HAVE ENTERED DEEPLY INTO THE INFESTED
STARPORT. BUT SOMETHING IS WRONG. THE
MONSTERS HAVE BROUGHT THEIR OWN REALITY
WITH THEM, AND THE STARPORT'S TECHNOLOGY
IS BEING SUBVERTED BY THEIR PRESENCE.

AHEAD, YOU SEE AN OUTPOST OF HELL, A
FORTIFIED ZONE. IF YOU CAN GET PAST IT,
YOU CAN PENETRATE INTO THE HAUNTED HEART
OF THE STARBASE AND FIND THE CONTROLLING
SWITCH WHICH HOLDS EARTH'S POPULATION
HOSTAGE. RROCK14 YOU HAVE WON! YOUR VICTORY HAS ENABLED
HUMANKIND TO EVACUATE EARTH AND ESCAPE
THE NIGHTMARE.  NOW YOU ARE THE ONLY
HUMAN LEFT ON THE FACE OF THE PLANET.
CANNIBAL MUTATIONS, CARNIVOROUS ALIENS,
AND EVIL SPIRITS ARE YOUR ONLY NEIGHBORS.
YOU SIT BACK AND WAIT FOR DEATH, CONTENT
THAT YOU HAVE SAVED YOUR SPECIES.

BUT THEN, EARTH CONTROL BEAMS DOWN A
MESSAGE FROM SPACE: "SENSORS HAVE LOCATED
THE SOURCE OF THE ALIEN INVASION. IF YOU
GO THERE, YOU MAY BE ABLE TO BLOCK THEIR
ENTRY.  THE ALIEN BASE IS IN THE HEART OF
YOUR OWN HOME CITY, NOT FAR FROM THE
STARPORT." SLOWLY AND PAINFULLY YOU GET
UP AND RETURN TO THE FRAY. RROCK07 YOU ARE AT THE CORRUPT HEART OF THE CITY,
SURROUNDED BY THE CORPSES OF YOUR ENEMIES.
YOU SEE NO WAY TO DESTROY THE CREATURES'
ENTRYWAY ON THIS SIDE, SO YOU CLENCH YOUR
TEETH AND PLUNGE THROUGH IT.

THERE MUST BE A WAY TO CLOSE IT ON THE
OTHER SIDE. WHAT DO YOU CARE IF YOU'VE
GOT TO GO THROUGH HELL TO GET TO IT? RROCK17 THE HORRENDOUS VISAGE OF THE BIGGEST
DEMON YOU'VE EVER SEEN CRUMBLES BEFORE
YOU, AFTER YOU PUMP YOUR ROCKETS INTO
HIS EXPOSED BRAIN. THE MONSTER SHRIVELS
UP AND DIES, ITS THRASHING LIMBS
DEVASTATING UNTOLD MILES OF HELL'S
SURFACE.

YOU'VE DONE IT. THE INVASION IS OVER.
EARTH IS SAVED. HELL IS A WRECK. YOU
WONDER WHERE BAD FOLKS WILL GO WHEN THEY
DIE, NOW. WIPING THE SWEAT FROM YOUR
FOREHEAD YOU BEGIN THE LONG TREK BACK
HOME. REBUILDING EARTH OUGHT TO BE A
LOT MORE FUN THAN RUINING IT WAS.
 RROCK13 CONGRATULATIONS, YOU'VE FOUND THE SECRET
LEVEL! LOOKS LIKE IT'S BEEN BUILT BY
HUMANS, RATHER THAN DEMONS. YOU WONDER
WHO THE INMATES OF THIS CORNER OF HELL
WILL BE. RROCK19 CONGRATULATIONS, YOU'VE FOUND THE
SUPER SECRET LEVEL!  YOU'D BETTER
BLAZE THROUGH THIS ONE!
 You've fought your way out of the infested
experimental labs.   It seems that UAC has
once again gulped it down.  With their
high turnover, it must be hard for poor
old UAC to buy corporate health insurance
nowadays..

Ahead lies the military complex, now
swarming with diseased horrors hot to get
their teeth into you. With luck, the
complex still has some warlike ordnance
laying around. You hear the grinding of heavy machinery
ahead.  You sure hope they're not stamping
out new hellspawn, but you're ready to
ream out a whole herd if you have to.
They might be planning a blood feast, but
you feel about as mean as two thousand
maniacs packed into one mad killer.

You don't plan to go down easy. The vista opening ahead looks real damn
familiar. Smells familiar, too -- like
fried excrement. You didn't like this
place before, and you sure as hell ain't
planning to like it now. The more you
brood on it, the madder you get.
Hefting your gun, an evil grin trickles
onto your face. Time to take some names. Suddenly, all is silent, from one horizon
to the other. The agonizing echo of Hell
fades away, the nightmare sky turns to
blue, the heaps of monster corpses start 
to evaporate along with the evil stench 
that filled the air. Jeeze, maybe you've
done it. Have you really won?

Something rumbles in the distance.
A blue light begins to glow inside the
ruined skull of the demon-spitter. What now? Looks totally different. Kind
of like King Tut's condo. Well,
whatever's here can't be any worse
than usual. Can it?  Or maybe it's best
to let sleeping gods lie.. Time for a vacation. You've burst the
bowels of hell and by golly you're ready
for a break. You mutter to yourself,
Maybe someone else can kick Hell's ass
next time around. Ahead lies a quiet town,
with peaceful flowing water, quaint
buildings, and presumably no Hellspawn.

As you step off the transport, you hear
the stomp of a cyberdemon's iron shoe. You gloat over the steaming carcass of the
Guardian.  With its death, you've wrested
the Accelerator from the stinking claws
of Hell.  You relax and glance around the
room.  Damn!  There was supposed to be at
least one working prototype, but you can't
see it. The demons must have taken it.

You must find the prototype, or all your
struggles will have been wasted. Keep
moving, keep fighting, keep killing.
Oh yes, keep living, too. Even the deadly Arch-Vile labyrinth could
not stop you, and you've gotten to the
prototype Accelerator which is soon
efficiently and permanently deactivated.

You're good at that kind of thing. You've bashed and battered your way into
the heart of the devil-hive.  Time for a
Search-and-Destroy mission, aimed at the
Gatekeeper, whose foul offspring is
cascading to Earth.  Yeah, he's bad. But
you know who's worse!

Grinning evilly, you check your gear, and
get ready to give the bastard a little Hell
of your own making! The Gatekeeper's evil face is splattered
all over the place.  As its tattered corpse
collapses, an inverted Gate forms and
sucks down the shards of the last
prototype Accelerator, not to mention the
few remaining demons.  You're done. Hell
has gone back to pounding bad dead folks 
instead of good live ones.  Remember to
tell your grandkids to put a rocket
launcher in your coffin. If you go to Hell
when you die, you'll need it for some
final cleaning-up ... You've found the second-hardest level we
got. Hope you have a saved game a level or
two previous.  If not, be prepared to die
aplenty. For master marines only. Betcha wondered just what WAS the hardest
level we had ready for ya?  Now you know.
No one gets out alive.       �T@     JS@     �S@     �U@     �S@     �T@     SKY2 SKY3 F_SKY1 Press escape to quit. G_CheckSpot: unexpected angle %d
 Only %i deathmatch spots, 4 required map31 wb recovery.dsg Failed to open either '%s' or '%s' to write savegame. Savegame buffer overrun Failed to open savegame file '%s' for writing.
But your game has been saved to '%s' for recovery. game saved. rb Bad savegame -maxdemo Doom 1.2 does not have a version code! v1.0/v1.1/v1.2 %i.%i (unknown) Demo is from a different game version!
(read %i, should be %i)

*** You may need to upgrade your version of Doom to v1.9. ***
    See: https://www.doomworld.com/classicdoom/info/patches.php
    This appears to be %s. -netdemo -nodraw timed %i gametics in %i realtics (%f fps) Demo %s recorded DOOM%02i.%s screen shot %s is turbo! consistency failure (%i should be %i) NET GAME SKY4 v1.4 v1.5 v1.6/v1.666 v1.7/v1.7a v1.8 v1.9         �v@     �v@     w@     w@     w@     w@     !w@     (w@     /w@             �B     �B     (�B                             -�B     2�B     7�B     C�B     N�B     S�B                                                                                                      �Qe     �Qe     �Qe     �Qe     |Qe     xQe     tQe     pQe       BSTCFN%.3d Unknown level [Message unsent] You mumble to yourself Who's there? You scare yourself You start to rave You've lost it... level 1: entryway level 2: underhalls level 3: the gantlet level 4: the focus level 5: the waste tunnels level 6: the crusher level 7: dead simple level 8: tricks and traps level 9: the pit level 10: refueling base level 11: 'o' of destruction! level 12: the factory level 13: downtown level 14: the inmost dens level 15: industrial zone level 16: suburbs level 17: tenements level 18: the courtyard level 19: the citadel level 20: gotcha! level 21: nirvana level 22: the catacombs level 23: barrels o' fun level 24: the chasm level 25: bloodfalls level 26: the abandoned mines level 27: monster condo level 28: the spirit world level 29: the living end level 30: icon of sin level 31: wolfenstein level 32: grosse level 1: congo level 2: well of souls level 3: aztec level 4: caged level 5: ghost town level 6: baron's lair level 7: caughtyard level 8: realm level 9: abattoire level 10: onslaught level 11: hunted level 12: speed level 13: the crypt level 14: genesis level 15: the twilight level 16: the omen level 17: compound level 18: neurosphere level 19: nme level 20: the death domain level 21: slayer level 22: impossible mission level 23: tombstone level 24: the final frontier level 25: the temple of darkness level 26: bunker level 27: anti-christ level 28: the sewers level 29: odyssey of noises level 30: the gateway of hell level 31: cyberden level 32: go 2 it level 1: system control level 2: human bbq level 3: power control level 4: wormhole level 5: hanger level 6: open season level 7: prison level 8: metal level 9: stronghold level 10: redemption level 11: storage facility level 12: crater level 13: nukage processing level 14: steel works level 15: dead zone level 16: deepest reaches level 17: processing area level 18: mill level 19: shipping/respawning level 20: central processing level 21: administration center level 22: habitat level 23: lunar mining project level 24: quarry level 25: baron's den level 26: ballistyx level 27: mount pain level 28: heck level 29: river styx level 30: last call level 31: pharaoh level 32: caribbean E1M1: Hangar E1M2: Nuclear Plant E1M3: Toxin Refinery E1M4: Command Control E1M5: Phobos Lab E1M6: Central Processing E1M7: Computer Station E1M8: Phobos Anomaly E1M9: Military Base E2M1: Deimos Anomaly E2M2: Containment Area E2M3: Refinery E2M4: Deimos Lab E2M5: Command Center E2M6: Halls of the Damned E2M7: Spawning Vats E2M8: Tower of Babel E2M9: Fortress of Mystery E3M1: Hell Keep E3M2: Slough of Despair E3M3: Pandemonium E3M4: House of Pain E3M5: Unholy Cathedral E3M6: Mt. Erebus E3M7: Limbo E3M8: Dis E3M9: Warrens E4M1: Hell Beneath E4M2: Perfect Hatred E4M3: Sever The Wicked E4M4: Unruly Evil E4M5: They Will Repent E4M6: Against Thee Wickedly E4M7: And Hell Followed E4M8: Unto The Cruel E4M9: Fear NEWLEVEL Green:  Indigo:  Brown:  Red:  No I'm ready to kick butt! I'm OK. I'm not looking too good! Help! You suck! Next time, scumbag... Come here! I'll take care of it. Yes TROO SHTG PUNG PISG PISF SHTF SHT2 CHGG CHGF MISG MISF SAWG PLSG PLSF BFGG BFGF BLUD PUFF BAL1 BAL2 PLSS PLSE MISL BFS1 BFE1 BFE2 TFOG IFOG PLAY POSS SPOS FIRE FATB FBXP SKEL MANF FATT CPOS SARG HEAD BAL7 BOSS BOS2 SKUL SPID BSPI APLS APBX CYBR PAIN SSWV KEEN BBRN BOSF ARM1 ARM2 BAR1 BEXP FCAN BON1 BON2 BKEY RKEY YKEY BSKU RSKU YSKU STIM MEDI PINV PSTR PINS MEGA SUIT PMAP PVIS CLIP AMMO BROK CELL CELP SHEL SBOX BPAK BFUG MGUN CSAW LAUN PLAS SHOT SGN2 COLU SMT2 GOR1 POL2 POL5 POL4 POL3 POL1 POL6 GOR2 GOR3 GOR4 GOR5 SMIT COL1 COL2 COL3 COL4 CAND CBRA COL6 TRE1 TRE2 ELEC CEYE FSKU COL5 TBLU TGRN TRED SMBT SMGT SMRT HDB1 HDB2 HDB3 HDB4 HDB5 HDB6 POB1 POB2 BRS1 TLMP TLP2 use_joystick joystick_index joystick_x_axis joystick_y_axis joystick_strafe_axis joystick_x_invert joystick_y_invert joystick_strafe_invert joystick_physical_button%i -nosound -nosfx -nomusic  Doom Generic is free software, covered by the GNU General Public
 License.  There is NO warranty; not even for MERCHANTABILITY or FITNESS
 FOR A PARTICULAR PURPOSE. You are welcome to change and distribute
 copies under certain conditions. See the source for more information. Warning: recursive call to I_Error detected.
 

 -nogui /usr/bin/zenity --help >/dev/null 2>&1 $`\! /usr/bin/zenity %s --error --text=%s -mb Unable to allocate %i MiB of RAM for zone zone memory: %p, %x allocated for zone
 -setmem dos622 dos71 dosbox     �           �� ep        W� �p  Unknown configuration variable: '%s' -config 	default file: %s
 saving config in %s
 -extraconfig         extra configuration file: %s
 Using %s for configuration and saves
 savegame/ Using %s for savegames
 graphical_startup autoadjust_video_settings fullscreen aspect_ratio_correct startup_delay screen_width screen_height screen_bpp grabmouse novert mouse_acceleration mouse_threshold snd_samplerate snd_cachesize snd_maxslicetime_ms snd_musiccmd opl_io_port png_screenshots vanilla_keyboard_mapping video_driver window_position joystick_physical_button0 joystick_physical_button1 joystick_physical_button2 joystick_physical_button3 joystick_physical_button4 joystick_physical_button5 joystick_physical_button6 joystick_physical_button7 joystick_physical_button8 joystick_physical_button9 joyb_strafeleft joyb_straferight joyb_menu_activate joyb_prevweapon joyb_nextweapon mouseb_strafeleft mouseb_straferight mouseb_use mouseb_backward mouseb_prevweapon mouseb_nextweapon dclick_use key_pause key_menu_activate key_menu_up key_menu_down key_menu_left key_menu_right key_menu_back key_menu_forward key_menu_confirm key_menu_abort key_menu_help key_menu_save key_menu_load key_menu_volume key_menu_detail key_menu_qsave key_menu_endgame key_menu_messages key_menu_qload key_menu_quit key_menu_gamma key_spy key_menu_incscreen key_menu_decscreen key_menu_screenshot key_map_toggle key_map_north key_map_south key_map_east key_map_west key_map_zoomin key_map_zoomout key_map_maxzoom key_map_follow key_map_grid key_map_mark key_map_clearmark key_weapon1 key_weapon2 key_weapon3 key_weapon4 key_weapon5 key_weapon6 key_weapon7 key_weapon8 key_prevweapon key_nextweapon key_arti_all key_arti_health key_arti_poisonbag key_arti_blastradius key_arti_teleport key_arti_teleportother key_arti_egg key_arti_invulnerability key_message_refresh key_demo_quit key_multi_msg key_multi_msgplayer1 key_multi_msgplayer2 key_multi_msgplayer3 key_multi_msgplayer4 key_multi_msgplayer5 key_multi_msgplayer6 key_multi_msgplayer7 key_multi_msgplayer8 show_talk voice_volume key_right key_left key_up key_down key_strafeleft key_straferight key_useHealth key_jump key_flyup key_flydown key_flycenter key_lookup key_lookdown key_lookcenter key_invquery key_mission key_invPop key_invKey key_invHome key_invEnd key_invleft key_invright key_invLeft key_invRight key_useartifact key_invUse key_invDrop key_lookUp key_lookDown key_fire key_use key_strafe key_speed use_mouse mouseb_fire mouseb_strafe mouseb_forward mouseb_jump joyb_fire joyb_strafe joyb_use joyb_speed joyb_jump screensize snd_musicdevice snd_sfxdevice snd_sbport snd_sbirq snd_sbdma snd_mport usegamma savedir messageson back_flat nickname chatmacro0 chatmacro1 chatmacro2 chatmacro3 chatmacro4 chatmacro5 chatmacro6 chatmacro7 chatmacro8 chatmacro9 comport                             #�@     #�@     �@     Y�@     3�@                                    1   2   3   4   5   6   7   8   9   0   -   =      	   q   w   e   r   t   y   u   i   o   p   [   ]      �   a   s   d   f   g   h   j   k   l   ;   '   `   �   \   z   x   c   v   b   n   m   ,   .   /   �   *   �       �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   -   �   5   �   +   �   �   �   �   �               �   �                                                                                                                                                       �       key_multi_msgplayer%i Messages OFF Messages ON HELP1 M_DOOM M_NEWG M_SKILL M_EPISOD empty slot HELP Unhandled game version High detail Low detail M_LSLEFT M_LSCNTR M_LSRGHT M_THERML M_THERMM M_THERMR M_THERMO M_SVOL M_OPTTTL M_CELL1 M_CELL2 you can't quickload during a netgame!

press a key. you haven't picked a quicksave slot yet!

press a key. do you want to quickload the game named

'%s'?

press y or n. you can't end a netgame!

press a key. are you sure you want to end the game?

press y or n. %s

(press y to quit to dos.) are you sure? this skill level
isn't even remotely fair.

press y or n. M_LOADG M_SAVEG _ you can't do load while in a net game!

press a key. you can't save if you aren't playing!

press a key. quicksave over your game named

'%s'?

press y or n. you can't start a new game
while in a network game.

press a key. this is the shareware version of doom.

you need to order the entire trilogy.

press a key. M_Episode: 4th episode requires UltimateDOOM
 M_MSGOFF M_MSGON M_GDHIGH M_GDLOW M_SKULL1 M_SKULL2    ��B     ��B     ��B     ��B     Couldn't read file %s  0x%x  0X%x  0%o Warning: Truncated '%s' lump name to '%.8s'.
 Failed to duplicate string (length %i)
 M_StringReplace: Failed to allocate new string M_StringJoin: Failed to allocate new string. /tmp                    m���kK���BJ�/P�̀�YM$_nU0Ԍ��O�2�4��xD�>F��[Ř��h���ʶ��Q��*'�����]z�� ��F�.��5�m���\��ME�N��Ԧq^�)2�1o�F<%�K��8*���I�M=bćj?��V`�qe���qP�l���Okp�g���x�:<R��B����QΣ-?Z�r;!�_�{b}�F��6m�G�]�W�4{�$.4��L�T%إ�j��b+'����Tv޻�x�����@     ��@     ��@     X�@     _�@     F�@     ��@     ��@     ��@     {�@     ]�@     {�@     ¿@     7�@     ¿@     ׿@     ׿@     �@     ׿@     �@     	�@     ��@     ��@     	�@     7�@     ��@     ��@     x�@     You need a blue key to activate this object You need a red key to activate this object You need a yellow key to activate this object You need a blue key to open this door You need a yellow key to open this door You need a red key to open this door EV_VerticalDoor: Tried to close something that wasn't a door.
 Weird actor->movedir! P_NewChaseDir: called with no target       ��@     ��@     �@     N�@     ��@     @�@     ��@     ��@     �@     F�@     ��@     d�@     ��@     P_GiveAmmo: bad type %i Picked up the armor. Picked up the MegaArmor! Picked up a health bonus. Picked up an armor bonus. Supercharge! MegaSphere! Picked up a blue keycard. Picked up a yellow keycard. Picked up a red keycard. Picked up a blue skull key. Picked up a yellow skull key. Picked up a red skull key. Picked up a stimpack. Picked up a medikit that you REALLY need! Picked up a medikit. Invulnerability! Berserk! Partial Invisibility Radiation Shielding Suit Computer Area Map Light Amplification Visor Picked up a clip. Picked up a box of bullets. Picked up a rocket. Picked up a box of rockets. Picked up an energy cell. Picked up an energy cell pack. Picked up 4 shotgun shells. Picked up a box of shotgun shells. Picked up a backpack full of ammo! You got the BFG9000!  Oh, yes. You got the chaingun! A chainsaw!  Find some meat! You got the rocket launcher! You got the plasma gun! You got the shotgun! You got the super shotgun! P_SpecialThing: Unknown gettable thing  q�@     ��@     �@     �@     �@     ��@     ��@     ��@     ��@     ��@     ��@     �@     �@     7�@     \�@     "�@     ��@     ��@     ��@     Q�@     �@      �@     >�@     Z�@     ��@     ��@     ��@     �@     1�@     [�@     ��@     ��@     ��@     �@     O�@     v�@     ��@     ��@     ��@     PTR_SlideTraverse: not a line? -spechit SpechitOverrun: Warning: unable to emulatean overrun where numspechit=%i
                                                                                                           �Vf                    �Jf                    �Jf                    �Jf                                    x                                                     0_f                                                                                  (        `f                                          l`f                                           H`f                    D`f                                           �`f                                     P_SpawnMapThing: Unknown type %i at (%i, %i) P_AddActivePlat: no more plats! P_RemoveActivePlat: can't find plat!       �,A     �,A     q,A     ),A     �,A     saveg_write8: Error while writing save game
 saveg_read8: Unexpected end of file while reading save game
 temp.dsg doomsav%d.dsg %s%s version %i P_UnarchiveSpecials:Unknown tclass %i in savegame      �MA     +NA     �NA     ,OA     �OA     KPA     �PA     ,QA     map0%i map%i PadRejectArray: REJECT lump too short to pad! (%i > %i)
 -reject_pad_with_ff P_CrossSubsector: ss %i with numss = %i P_InitPicAnims: bad cycle from %s to %s Sector with more than 22 adjoining sectors. Vanilla will crash here P_PlayerInSpecialSector: unknown special %i EV_DoDonut: linedef had no second sidedef! Unexpected behavior may occur in Vanilla Doom. 
 EV_DoDonut: WARNING: emulating buffer overrun due to NULL back sector. Unexpected behavior may occur in Vanilla Doom.
 -donut DonutOverrun: The second parameter for "-donut" switch should be greater than 0 and less than number of flats (%d). Using default value (%d) instead. 
 Too many scrolling wall linedefs! (Vanilla limit is 64)     EfA     LfA     ^fA     bfA     lfA     �hA     vfA     �hA     }fA     �hA     �fA     �fA     �hA     �hA     �fA     �fA     �hA     �fA     �hA     �hA     �fA     �hA     �hA     �fA     �hA     �hA     �hA     �hA     �fA     �hA     �hA     �hA     �hA     �fA     �fA     �fA     gA     �gA     �fA     �hA     �hA     �hA     gA     �hA     �hA     �hA     �hA     �hA     �hA     �hA     gA     gA     "gA     �hA     /gA     9gA     FgA     MgA     �hA     �hA     �hA     �hA     �hA     �hA     �hA     �hA     �hA     �hA     �hA     �hA     �gA     �gA     �gA     hA     hA     hA     �hA     hA     $hA     /hA     6hA     @hA     GhA     �hA     QhA     XhA     ^hA     ghA     phA     thA     {hA     �hA     �hA     �hA     �hA     �hA     �hA     �hA     rgA     �hA     �hA     �hA     TgA     �hA     �hA     �hA     ^gA     hgA     �gA     �hA     �hA     �hA     �hA     �hA     �hA     �hA     �hA     �gA     �hA     �gA     �hA     �hA     �gA     �gA     �hA     �hA     �hA     �hA     �gA     �hA     �hA     �hA     �hA     �hA     �hA     �hA     �hA     �hA     �hA     �gA     �iA     �iA     0jA     �iA     0jA     �iA     0jA     jA     0jA     0jA     0jA     0jA     �iA     2nA     <nA     @nA     QnA     �nA     �nA     �nA     hnA     rnA     znA     �nA     �nA     �nA     �nA     �nA     �nA     �nA     P_StartButton: no button slots left!    ?rA     wtA     wtA     wtA     wtA     wtA     OrA     wtA     hrA     wtA     rrA     wtA     wtA     �rA     �rA     wtA     wtA     �rA     wtA     �rA     �rA     wtA     �rA     wtA     wtA     ?rA     ?rA     ?rA     �rA     wtA     ?rA     ?rA     ?rA     ?rA     wtA     wtA     wtA     wtA     wtA     wtA     �rA     zsA     �sA     wtA     �sA     wtA     wtA     wtA     �rA     �rA     �rA     wtA     wtA     wtA     sA     wtA     wtA     wtA     wtA     �sA     �sA     �sA     �sA     �sA     �sA     �sA     �sA     �sA     �sA     �sA     �rA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     DtA     wtA     sA     sA     sA     wtA     wtA     wtA     wtA     wtA     wtA     wtA     sA     %sA     ,sA      tA     
tA     tA     ?rA     ?rA     wtA     wtA     wtA     >sA     tA     wtA     wtA     wtA     JsA     wtA     wtA     wtA     TsA     2tA     ^sA     DtA     ^sA     DtA     ^sA     VtA     ]tA     psA     R_Subsector: ss %i with numss = %i r_data.c R_GenerateLookup: column without a patch (%s)
 R_GenerateLookup: texture %i is >64k PNAMES TEXTURE1 TEXTURE2 S_END R_InitTextures: bad texture directory R_InitTextures: Missing patch in texture %s F_START COLORMAP R_FlatNumForName: %s not found R_TextureNumForName: %s not found R_DrawColumn: %i to %i at %i R_DrawFuzzColumn: %i to %i at %i R_DrawSpan: %i to %i at %i GRNROCK FLOOR7_2 brdr_t brdr_b brdr_l brdr_r brdr_tl brdr_tr brdr_bl brdr_br R_MapPlane: %i, %i at %i R_FindPlane: no more visplanes R_DrawPlanes: drawsegs overflow (%i) R_DrawPlanes: visplane overflow (%i) R_DrawPlanes: opening overflow (%i) Bad R_RenderWallRange: %i to %i R_InstallSpriteLump: Bad frame characters in lump %i R_InitSprites: Sprite %s frame %c has multip rot=0 lump R_InitSprites: Sprite %s frame %c has rotations and a rot=0 lump R_InitSprites: Sprite %s : %c : %c has two lumps mapped to it R_InitSprites: No patches found for %s frame %c R_InitSprites: Sprite %s frame %c is missing rotations R_DrawSpriteRange: bad texturecolumn R_ProjectSprite: invalid sprite number %i  R_ProjectSprite: invalid sprite frame %i : %i  e1m1 e1m2 e1m3 e1m4 e1m5 e1m6 e1m7 e1m8 e1m9 e2m1 e2m2 e2m3 e2m4 e2m5 e2m6 e2m7 e2m8 e2m9 e3m1 e3m2 e3m3 e3m4 e3m5 e3m6 e3m7 e3m8 e3m9 inter intro bunny victor introa runnin stalks countd betwee the_da shawn ddtblu in_cit dead stlks2 theda2 ddtbl2 runni2 dead2 stlks3 romero shawn2 messag count2 ddtbl3 ampie theda3 adrian messg2 romer2 tense shawn3 openin evil ultima read_m dm2ttl dm2int STTMINUS drawNum: n->y - ST_Y < 0 updateMultIcon: y - ST_Y < 0 updateBinIcon: y - ST_Y < 0 STTNUM%d STYSNUM%d STTPRCNT STKEYS%d STARMS STGNUM%d STFB%d STBAR STFST%d%d STFTR%d0 STFTL%d0 STFOUCH%d STFEVL%d STFKILL%d STFGOD0 STFDEAD0 Degreelessness Mode On Degreelessness Mode Off Ammo (no keys) Added Very Happy Ammo Added Music Change IMPOSSIBLE SELECTION No Clipping Mode ON No Clipping Mode OFF Power-up Toggled inVuln, Str, Inviso, Rad, Allmap, or Lite-amp ... doesn't suck - GM ang=0x%x;x,y=(0x%x,0x%x) Changing Level... Bad sfx #: %d Attempt to set music volume at %d Attempt to set sfx volume at %d Bad music number %d d_%s                                             	                               	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������
 !"$%&'()*,-./012346789:;<=>?@ABCEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������	 !#$&'(*+-./02346789;<=>?ABCDEFHIJKLMNOPRSTUVWXYZ[\]^_`abdefghijklmnopqrrstuvwxyz{|}~�����������������������������������������������������������������������������������������������������������������������������������������������������������"$&()+-/124579:<=?@ACDFGHJKLMOPQRTUVWXZ[\]^_`bcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������� $'*-02579<>@BDEGIKLNPQSTVWYZ\]^`abdefgijklmnpqrstuvwxyz{|}~�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������    � �/
 cG ._ �v  ��# S�( �- ��2 �8 c= #5B �LG �dL U|Q �V ��[ p�` �e ��j p
p "u �9z PQ �h� }�� �� ��� ǘ �ޝ �� �� 	%� w<� �S� Ak� ��� �� C�� ��� ��� �� B� p%� �<� �S� �j� �� �� ��������v"D9"
P'�f,x}1 �6��;V�@��Eb�J�PFU�1Z H_L^d�tin�s�x�}&� ����$��:��P�Nf��{����4�����4Һ�����N��'��<��Q��f�|������������B�����"�6�JL_�s ̇%��*�/�4��9��>��CdI'N�:S,NX�a] ubL�g��l��q��v��{�����D����2�E��W��i�(|�\��x�����tĽP�������d���T.��?��P�b�$s� ����̥����	���`���#�((�8-�H2HX7�g<twA�F<�Kx�P��U��Z��_d�d�i��n<t�y�)~8�0F�(T� b��o�d}�슡T�����в�俵�̺�ٿl���������,�T$�X0�@<�H��S�<_��j��u �0����� ���$��) �.�3��8��=h�B�HPM�R�"W�+\�4a@=f�EkHNp�Vu�^z�f�n��v� ~�������0��@��(��������p�����������h���������� ����������8�����
 �� X �%�"*x%/0(4�*9(->h/C�1Hp3M05R�6W@8\�9a�:f�;k`<p =up=z�=�=��=��=�@=��<��;�;�:��8�h7��5�4�(2�0��-�`+��(��%� #������X�x�p�8	�8 x���`����#��(�-��2��7P�<��A�F�K��PX�UȝZ�_�d��i�}n ushlx�c}hZ�Q��G��=�4��)���8��
�������P��ݽ(��H��8����p�����؇��z�xm��_�8R�PD�06��'H�
��`� �h� ��%��*X�/�48|9Xk>@ZC�HHp7M�%R�W�\0�`��e��j��op�t��y@|~Ph�0T��?�8+�h�X���֥����Ȕ�`~��g��P��9��"� �8��8�� �����ؑ��x��_�`F��,�������� � ��r PW%�;*�/`4��80�=@�B�G�rL UQ7V�[��_��d �i��n�~s�^x ?}������݋����z� Y� 7����в@�� ���f� C�@� ����� ��@�� h��B�� ��������Ѓ 	�\	�5
	0	��	��	@�	�m"	�D'	�,	��0	�5	0�:	 u?	�JD	  I	@�M	�R	��W	 s\	 Ga	�f	P�j	��o	��t	0gy	�9~	��	�݇	@��	���	�Q�	p"�	 �	@ä	0��	�b�	P2�	��	Pм	��	@m�	P;�		�	���	���	�p�	P=�	�	�	���	���	 m�	`8�	P 
 �
`�	
�b
P,
��
 �
 �!
�P&
@+
P�/
0�4
�p9
 8>
��B
��G
 �L
 RQ
�V
��Z
��_
�gd
P,i
��m
��r
�xw
 <|
0��
 
���
 G�
 	�
�ʘ
0��
PM�
 �
�Ϋ
���
�N�
��
�;
���
�K�

�
@��
��
�C�
� �
н�
�z�
�6�
���
���
 j�
 % ���
�T�@����:"0�&��+�c0p5��9 �>�@C`�G��L�cQ V`�Z`�_ 8d`�hp�m Tr�w��{pm���҉���p5������ H�`��P���W�@�@���d�P�P��o�p����@v��"�����z�&�@��|��&�����z $P�0v����np$��(�d-02��6pW;�?P�D@GI��M0�R04W��[ {`e��icn s��w H|������)��Ɏ�i���ড়�F������` �����Z�P������/� ��pf�`���06� ���i���Л�`4�����d� �0�*���V�� � "�&`@+p�/0h4��8��=`!B��F�EKp�O�hT��Xp�]�b��f@:kp�o`Xt��xu}��p����P���6���N� ڡ e��� z� ���������P(����`8��� G����0T�P�� `�`��`j� ��@s�0� �z �	ЀPp�@�� �	%`�)�
.��2P
7��;p@��D I��M` Rp}V0�Z�v_��c nh`�l@dq��u Yz��~0L�PŇ >�P��P.�ख़ � ���
����p���k����U�����=�P���$�P���	��{�����^����p@����� � �� ���m@�0Jз%�p��j#P�'�A,��0`5��9��= UB �F�&K@�O@�S�^X �\ -a��e��iP_n��r�)wP�{��`V�й����� ��C�������g��ǫ (���� ��E�p����P`������Pw����p/���� ���@� ������N����� �X���_�� @c!�%@* c.��2�7�_; �? D�XH�L��P@NU@�Y �]@@b �f��j�.o�}s��w�|`g����`��M����`��0�`{��Ţ���Y�ࢯ��@4�`|� ��`�@R���� ���$� j� ������7��{������D������  
 K	����� K ���" ' E+`�/��3 �7`8<`t@��D��H�%M�_Q��U@�Y`^ Eb`}f@�j��n $s�Zw �{��`���1�@f�����Δ � 5��g�@�� ̩����.��_����࿾`����@M��{���� �� ��0� ]� ���������
��4��^�@�`� �	`@*�Q�x����"��& +@6/ [3@7 �;��?��C@H�.L`PP�qT��X��\��`��d i 2m�Pq�nu��y �} ǁ������� 7� R��l����`������Ҫ@�`� �`2�@I��_��u��������� ��@����� � �`*�`<� N�@_� p�`� `� � ��@� ����� �%�)�-@%1@05 ;9@E= OA�XE�aI jM`rQ zU��Y��] �a@�e �i`�m`�q�u �y��} ��ළ`��`�� ��`�� ��������@��`��@�������� ��@�� ��@�� ��������`�������� �� ���z��r��j� b� Y��O��E`;�0	�% @�@� � ��$��( �,`�0 �4��8��< p@ _D�MH@<L *P�T�X`�[��_��c�g��k��o�ts�^w�G{�0`���@��Ў`����� ���i��N��3� � ���߱�µ��� ���i�`K��,�@����`���������j��H��&������`�����@u��P��+  �
�� ��k@D`��! �%�)@x- N1�#5��8��<�@�uD IH@L��O �S��W`d[@5_�c �f��j un Dr�v��y@�}�{�`H����������w��B����֟`���i� 2����`²����P��������� i� .��������z��=�� �@��`�� G�`�@������I�`	���`��E	�@�`~ ;��`��n# *'��*��.�X2 6 �9��= <A��D �H bL�P��S��W�9[��^ �b@Wf�
j �m qq`#u`�x �| 8���@��@I����৒�V������@`�@� �� f� �`��`h� �@�� g�`�@���a��	�����X����@��`L� ��@�� <������� (�`�� n �`� T ��� 6 ��u�!@�$�Q(`�+��/�)3��6�b:��=��A�4E��H�iL`P��S�5W �Z@f^ �a@�e ,i��l�Xp`�s��w�{�~�@��ԅ�g�������������A�`Ҟ�b��� ��@� ��@.�@���I��־�c�����{� � �������0� �� C�����S���� c� ���p�����|����@	`� ��`�� ��!� %��(@",@�/ "3@�6  :��=�A �D`H@�K�O��R@V`�Y@�\�x`��c lg`�j ^n��q�Nu �x =|�@*�@�����������s���`[��Ξ@A����`%���� ��x� ��X�`Ƚ�7�@����`����� ]�����5����@�`x� ��@M� ��� ����`���Z�����) ����]��@)@���@W � �$��'@�*�F.`�1�	5�j8��;�+?��B �E@JI�L P eS��V�Z@|]��``4d��g �j�En �q��t`Sx��{ �]�`���� d���� � g������`f������@b�`�� ��Z�`�� �� O� ��`��`@���� �� .�`|�`�� �@e� ������J�@�����`,��v�����
��S ��@�`-
 u`�`�I ��� ! `$��'��*�,. p1 �4��7 8;�y>@�A`�D =H@}K@�N��Q�;U�zX�[��^`4b�qe@�h��k�&o@br��u@�x�|�L`�������� 1� i�ࠒ@ؕ ��E��{���� � ��P�������@�@� R�@�� ��������I� z���������7� f� ����� ����`H��t�@��������@!��K@u��������@@h`� ���!�% ((`M+ r.��1��4`�7�;�$>@GA`iD@�G��J��M`�P�T�.W NZ m]��`@�c@�f��i m  p�<s�Xv@ty��|�� ł`߅@�����+�`D��\��t�@��`�� ���Ф��`�����&� ;�@O� c��v���� ��`��`����� �����@�@��#�@3� B��P��^��l� z� ����� ��������� `�����	������`�`��$"�+% 2(�7+�=.�B1�G4 L7 P:�S=@W@@ZC�\F _I aL�bO�cR�dU�dX�d[�d^�ca�bd`ag�_j`]m�Zp�Ws�Tv Qy M|�H�C��>�@9�`3�@-��&���`�����@ ����`����ګ�Ю Ʊ ����� �� ������~��q� d�@V� H�`9�`*� �`�`����� �� ��������`������m��Z��F��2�`�	`� �	 ��@�`� n�V`> &!`$@�&��) �,�/@�2`q5 V8�:;�>`A��C��F@�I��L`oO�PR 2U�X`�Z��]@�`��c�qf`Pi�.l�o`�q��t��w �z@]} 9������ʈ �� ��X� 2� ��� �� ���k� C���`��ƭ`���q� G���@�`ľ ���k��>� ������� ��`X�@)���� �� ���i��8��� �� ���q�@?�`� ������q�@=���@�
�h�2 �`�@��V �� ��#�u&�<) , �.��1`T4�7@�9��<�f?�*B��D�G�sJ 6M �O��R {U <X��Z�]�|`�<c��e��h@yk�7n`�p �s pv -y��{��~�a� �@؆ ���M������ {�@4� �`���]�`��̤����:� � ���\�@�`Ƿ |��0���@���K����`���c�������x��)��������:���� �� I���� �� T��� �� \��� �� a � � c� � b� � ^� � W ��" �%@M(��*@�-@@0 �2`�5`08 �:`y=�@ �B�dE�H`�J�LM��O��R 2U �W�sZ@]`�_ Tb��d��g`1j��l no�r@�t�Fw@�y�| ���@S���`���#� �� X�������#�`���T��� ������� I�`߭`u� �����5�@ʺ�^���`�������?� ��@d� ���������� :�`��@Z���� y� �����$����@�����Z���� t�                                   K   }   �   �     F  x  �  �    B  t  �  �    =  o  �  �    8  j  �  �    3  f  �  �  �  /  a  �  �  �  *  \  �  �  �  %  W  �  �  �   	  S	  �	  �	  �	  
  N
  �
  �
  �
    I  {  �  �    D  v  �  �    ?  q  �  �    :  l  �  �    5  g  �  �  �  0  b  �  �  �  *  ]  �  �  �  %  W  �  �  �     R  �  �  �    M    �  �    G  y  �  �    A  t  �  �  
  <  n  �  �    6  h  �  �  �  0  b  �  �  �  *  \  �  �  �  $  V  �  �  �    P  �  �  �    J  |  �  �    C  u  �  �    =  o  �  �     6   h   �   �   �   0!  a!  �!  �!  �!  )"  Z"  �"  �"  �"  "#  S#  �#  �#  �#  $  L$  ~$  �$  �$  %  E%  w%  �%  �%  &  >&  o&  �&  �&  '  6'  h'  �'  �'  �'  .(  `(  �(  �(  �(  &)  X)  �)  �)  �)  *  P*  �*  �*  �*  +  H+  y+  �+  �+  ,  ?,  q,  �,  �,  -  7-  h-  �-  �-  �-  ..  `.  �.  �.  �.  %/  W/  �/  �/  �/  0  N0  0  �0  �0  1  D1  v1  �1  �1  
2  ;2  l2  �2  �2   3  13  b3  �3  �3  �3  '4  Y4  �4  �4  �4  5  O5  �5  �5  �5  6  D6  u6  �6  �6  	7  :7  k7  �7  �7  �7  /8  `8  �8  �8  �8  $9  U9  �9  �9  �9  :  J:  {:  �:  �:  ;  ?;  o;  �;  �;  <  3<  d<  �<  �<  �<  '=  X=  �=  �=  �=  >  L>  }>  �>  �>  ?  ??  p?  �?  �?  @  3@  d@  �@  �@  �@  &A  WA  �A  �A  �A  B  JB  zB  �B  �B  C  <C  mC  �C  �C  �C  /D  _D  �D  �D  �D  !E  QE  �E  �E  �E  F  CF  sF  �F  �F  G  4G  eG  �G  �G  �G  &H  VH  �H  �H  �H  I  GI  wI  �I  �I  J  8J  hJ  �J  �J  �J  (K  XK  �K  �K  �K  L  HL  xL  �L  �L  M  8M  hM  �M  �M  �M  'N  WN  �N  �N  �N  O  FO  vO  �O  �O  P  5P  eP  �P  �P  �P  $Q  SQ  �Q  �Q  �Q  R  AR  qR  �R  �R   S  /S  _S  �S  �S  �S  T  LT  |T  �T  �T  
U  9U  iU  �U  �U  �U  &V  VV  �V  �V  �V  W  BW  qW  �W  �W  �W  .X  ]X  �X  �X  �X  Y  IY  xY  �Y  �Y  Z  4Z  cZ  �Z  �Z  �Z  [  N[  }[  �[  �[  
\  9\  h\  �\  �\  �\  #]  R]  �]  �]  �]  ^  <^  k^  �^  �^  �^  %_  T_  �_  �_  �_  `  =`  l`  �`  �`  �`  &a  Ta  �a  �a  �a  b  =b  kb  �b  �b  �b  %c  Sc  �c  �c  �c  d  :d  id  �d  �d  �d  !e  Pe  ~e  �e  �e  f  6f  df  �f  �f  �f  g  Jg  xg  �g  �g  h  0h  ^h  �h  �h  �h  i  Ci  qi  �i  �i  �i  (j  Vj  �j  �j  �j  k  :k  hk  �k  �k  �k  l  Ll  zl  �l  �l  m  0m  ]m  �m  �m  �m  n  @n  mn  �n  �n  �n  #o  Po  }o  �o  �o  p  2p  _p  �p  �p  �p  q  Aq  nq  �q  �q  �q  "r  Or  |r  �r  �r  s  0s  ]s  �s  �s  �s  t  =t  it  �t  �t  �t  u  Iu  vu  �u  �u  �u  (v  Uv  �v  �v  �v  w  3w  `w  �w  �w  �w  x  >x  jx  �x  �x  �x  y  Hy  ty  �y  �y  �y  %z  Qz  }z  �z  �z  {  .{  Z{  �{  �{  �{  
|  6|  b|  �|  �|  �|  }  =}  i}  �}  �}  �}  ~  D~  p~  �~  �~  �~    J  v  �  �  �  $�  O�  {�  ��  Ҁ  ��  )�  T�  �  ��  ց  �  -�  X�  ��  ��  ڂ  �  0�  [�  ��  ��  ܃  �  3�  ^�  ��  ��  ߄  	�  4�  _�  ��  ��  ��  �  6�  `�  ��  ��  �  �  6�  a�  ��  ��  �  �  6�  `�  ��  ��  ��  
�  5�  _�  ��  ��  މ  	�  3�  ]�  ��  ��  ܊  �  1�  [�  ��  ��  ً  �  -�  W�  ��  ��  Ռ  ��  )�  S�  }�  ��  э  ��  $�  N�  x�  ��  ˎ  ��  �  I�  r�  ��  ŏ  �  �  B�  l�  ��  ��  �  �  ;�  d�  ��  ��  ��  
�  3�  \�  ��  ��  ؒ  �  *�  S�  |�  ��  Γ  ��   �  I�  r�  ��  Ĕ  �  �  ?�  h�  ��  ��  �  �  3�  \�  ��  ��  ֖  ��  '�  P�  x�  ��  ɗ  �  �  C�  k�  ��  ��  �  �  5�  ]�  ��  ��  ֙  ��  &�  N�  v�  ��  ƚ  �  �  >�  f�  ��  ��  ޛ  �  .�  U�  }�  ��  ͜  ��  �  D�  l�  ��  ��  �  
�  1�  Y�  ��  ��  Ϟ  ��  �  E�  m�  ��  ��  �  
�  1�  X�  �  ��  Π  ��  �  C�  j�  ��  ��  ߡ  �  -�  T�  {�  ��  Ȣ  �  �  <�  c�  ��  ��  ף  ��  $�  K�  q�  ��  ��  �  �  2�  X�  ~�  ��  ˥  �  �  >�  d�  ��  ��  צ  ��  #�  I�  o�  ��  ��  �  �  -�  S�  x�  ��  Ĩ  �  �  5�  [�  ��  ��  ̩  �  �  =�  b�  ��  ��  Ӫ  ��  �  C�  h�  ��  ��  ث  ��  #�  H�  m�  ��  ��  ܬ  �  &�  K�  p�  ��  ��  ߭  �  )�  N�  s�  ��  ��  �  �  *�  O�  s�  ��  ��  �  �  *�  O�  s�  ��  ��  �  �  )�  M�  q�  ��  ��  ޱ  �  &�  J�  n�  ��  ��  ڲ  ��  "�  F�  j�  ��  ��  ճ  ��  �  A�  d�  ��  ��  ϴ  �  �  :�  ]�  ��  ��  ȵ  �  �  2�  U�  x�  ��  ��  �  �  (�  K�  n�  ��  ��  ׷  ��  �  @�  c�  ��  ��  ̸  �  �  4�  V�  y�  ��  ��  �  �  &�  H�  k�  ��  ��  Һ  ��  �  9�  [�  ~�  ��  »  �  �  (�  J�  m�  ��  ��  Ҽ  ��  �  8�  Z�  |�  ��  ��  �  �  $�  F�  h�  ��  ��  ̾  �  �  1�  R�  t�  ��  ��  ؿ  ��  �  ;�  \�  ~�  ��  ��  ��  �  #�  D�  e�  ��  ��  ��  ��  	�  *�  K�  k�  ��  ��  ��  ��  �  /�  P�  p�  ��  ��  ��  ��  �  2�  S�  s�  ��  ��  ��  ��  �  4�  T�  t�  ��  ��  ��  ��  �  3�  S�  s�  ��  ��  ��  ��  �  1�  P�  p�  ��  ��  ��  ��  �  ,�  L�  k�  ��  ��  ��  ��  �  &�  E�  d�  ��  ��  ��  ��  ��  �  =�  [�  z�  ��  ��  ��  ��  �  2�  Q�  o�  ��  ��  ��  ��  �  &�  D�  b�  ��  ��  ��  ��  ��  �  6�  T�  r�  ��  ��  ��  ��  �  %�  C�  `�  ~�  ��  ��  ��  ��  �  0�  M�  k�  ��  ��  ��  ��  ��  �  8�  V�  s�  ��  ��  ��  ��  �  !�  >�  [�  x�  ��  ��  ��  ��  �  %�  B�  ^�  {�  ��  ��  ��  ��  
�  &�  B�  _�  {�  ��  ��  ��  ��  �  $�  A�  ]�  y�  ��  ��  ��  ��  �   �  <�  X�  t�  ��  ��  ��  ��  ��  �  5�  Q�  l�  ��  ��  ��  ��  ��  �  ,�  G�  b�  }�  ��  ��  ��  ��  �  �  :�  U�  p�  ��  ��  ��  ��  ��  �  +�  F�  `�  {�  ��  ��  ��  ��  ��  �  4�  N�  h�  ��  ��  ��  ��  ��  �  �  9�  S�  m�  ��  ��  ��  ��  ��  �  !�  ;�  T�  n�  ��  ��  ��  ��  ��  �   �  9�  S�  l�  ��  ��  ��  ��  ��  �  �  5�  N�  g�  �  ��  ��  ��  ��  ��  �  -�  E�  ^�  v�  ��  ��  ��  ��  ��  	�  !�  :�  R�  j�  ��  ��  ��  ��  ��  ��  �  *�  B�  Z�  r�  ��  ��  ��  ��  ��   �  �  /�  G�  ^�  v�  ��  ��  ��  ��  ��  �  �  0�  G�  _�  v�  ��  ��  ��  ��  ��  ��  �  -�  D�  [�  q�  ��  ��  ��  ��  ��  ��  �  &�  <�  R�  i�  �  ��  ��  ��  ��  ��  �  �  0�  F�  \�  r�  ��  ��  ��  ��  ��  ��  
�   �  6�  K�  a�  v�  ��  ��  ��  ��  ��  ��  �  !�  6�  K�  `�  u�  ��  ��  ��  ��  ��  ��  �  �  1�  F�  [�  o�  ��  ��  ��  ��  ��  ��  ��  �  (�  <�  P�  d�  y�  ��  ��  ��  ��  ��  ��  �  �  -�  A�  T�  h�  |�  ��  ��  ��  ��  ��  ��  �  �  ,�  ?�  S�  f�  y�  ��  ��  ��  ��  ��  ��  ��  �  %�  8�  K�  ^�  q�  ��  ��  ��  ��  ��  ��  ��  �  �  +�  =�  O�  b�  t�  ��  ��  ��  ��  ��  ��  ��  �  �  )�  ;�  M�  _�  q�  ��  ��  ��  ��  ��  ��  ��  ��  �  !�  2�  C�  U�  f�  w�  ��  ��  ��  ��  ��  ��  ��   �  �  "�  3�  D�  T�  e�  v�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  +�  <�  L�  \�  l�  |�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  +�  ;�  K�  Z�  j�  y�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  "�  1�  @�  O�  ^�  m�  |�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  ,�  ;�  I�  X�  f�  t�  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  +�  8�  F�  T�  b�  o�  }�  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  *�  7�  D�  Q�  ^�  k�  x�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  (�  5�  A�  M�  Z�  f�  r�  ~�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  #�  /�  ;�  F�  Q�  ]�  h�  s�  �  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  #�  .�  9�  C�  N�  X�  c�  m�  x�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  #�  -�  6�  @�  J�  S�  ]�  f�  p�  y�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  �  %�  .�  6�  ?�  H�  P�  Y�  a�  i�  r�  z�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  	�  �  �   �  (�  /�  6�  >�  E�  L�  T�  [�  b�  i�  p�  w�  �  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  	�  �  �  �  "�  (�  .�  4�  :�  @�  F�  K�  Q�  W�  ]�  b�  h�  m�  s�  x�  ~�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  �  �  �  �  !�  %�  )�  -�  1�  5�  9�  =�  A�  E�  H�  L�  P�  S�  W�  [�  ^�  b�  e�  i�  l�  o�  s�  v�  y�  |�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  |�  y�  v�  s�  o�  l�  i�  e�  b�  ^�  [�  W�  S�  P�  L�  H�  E�  A�  =�  9�  5�  1�  -�  )�  %�  !�  �  �  �  �  �  �  �  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ~�  x�  s�  m�  h�  b�  ]�  W�  Q�  K�  F�  @�  :�  4�  .�  (�  "�  �  �  �  	�  �  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  w�  p�  i�  b�  [�  T�  L�  E�  >�  6�  /�  (�   �  �  �  	�  �  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  z�  r�  i�  a�  X�  P�  H�  ?�  6�  .�  %�  �  �  �  �  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  y�  p�  f�  ]�  S�  J�  @�  6�  -�  #�  �  �  �  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  x�  m�  c�  X�  N�  C�  9�  .�  #�  �  �  �  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  s�  h�  ]�  Q�  F�  ;�  /�  #�  �  �  �  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ~�  r�  f�  Z�  M�  A�  5�  (�  �  �  �  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  x�  k�  ^�  Q�  D�  7�  *�  �  �  �  ��  ��  ��  ��  ��  ��  ��  ��  ��  }�  o�  b�  T�  F�  8�  +�  �  �  �  ��  ��  ��  ��  ��  ��  ��  ��  ��  t�  f�  X�  I�  ;�  ,�  �  �  �  ��  ��  ��  ��  ��  ��  ��  ��  |�  m�  ^�  O�  @�  1�  "�  �  �  ��  ��  ��  ��  ��  ��  ��  ��  y�  j�  Z�  K�  ;�  +�  �  �  ��  ��  ��  ��  ��  ��  ��  ��  |�  l�  \�  L�  <�  +�  �  �  ��  ��  ��  ��  ��  ��  ��  ��  v�  e�  T�  D�  3�  "�  �   �  ��  ��  ��  ��  ��  ��  ��  w�  f�  U�  C�  2�  !�  �  ��  ��  ��  ��  ��  ��  ��  ��  q�  _�  M�  ;�  )�  �  �  ��  ��  ��  ��  ��  ��  ��  t�  b�  O�  =�  +�  �  �  ��  ��  ��  ��  ��  ��  ��  q�  ^�  K�  8�  %�  �  ��  ��  ��  ��  ��  ��  ��  y�  f�  S�  ?�  ,�  �  �  ��  ��  ��  ��  ��  ��  |�  h�  T�  A�  -�  �  �  ��  ��  ��  ��  ��  ��  y�  d�  P�  <�  (�  �  ��  ��  ��  ��  ��  ��  ��  o�  [�  F�  1�  �  �  ��  ��  ��  ��  ��  ��  u�  `�  K�  6�  !�  �  ��  ��  ��  ��  ��  ��  v�  a�  K�  6�   �  
�  ��  ��  ��  ��  ��  ��  r�  \�  F�  0�  �  �  ��  ��  ��  ��  ��  �  i�  R�  <�  &�  �  ��  ��  ��  ��  ��  ��  q�  [�  D�  -�  �  ��  ��  ��  ��  ��  ��  v�  _�  G�  0�  �  �  ��  ��  ��  ��  ��  v�  ^�  G�  /�  �   �  ��  ��  ��  ��  ��  r�  Z�  B�  *�  �  ��  ��  ��  ��  ��  ��  j�  R�  :�  !�  	�  ��  ��  ��  ��  ��  v�  ^�  E�  -�  �  ��  ��  ��  ��  ��  �  g�  N�  5�  �  �  ��  ��  ��  ��  ��  l�  S�  9�   �  �  ��  ��  ��  ��  ��  n�  T�  ;�  !�  �  ��  ��  ��  ��  ��  m�  S�  9�  �  �  ��  ��  ��  ��  ��  h�  N�  4�  �  ��  ��  ��  ��  ��  {�  `�  F�  +�  �  ��  ��  ��  ��  ��  p�  U�  :�  �  �  ��  ��  ��  ��  }�  b�  G�  ,�  �  ��  ��  ��  ��  ��  l�  Q�  5�  �  ��  ��  ��  ��  ��  t�  X�  <�   �  �  ��  ��  ��  ��  y�  ]�  A�  $�  �  ��  ��  ��  ��  {�  _�  B�  &�  
�  ��  ��  ��  ��  {�  ^�  B�  %�  �  ��  ��  ��  ��  x�  [�  >�  !�  �  ��  ��  ��  ��  s�  V�  8�  �  ��  ��  ��  ��  ��  k�  M�  0�  �  ��  ��  ��  ��  ~�  `�  C�  %�  �  ��  ��  ��  ��  r�  T�  6�  �  ��  ��  ��  ��  ��  b�  D�  &�  �  ��  ��  ��  ��  o�  Q�  2�  �  ��  ��  ��  ��  z�  [�  =�  �  ��  ��  ��  ��  ��  d�  E�  &�  �  ��  ��  ��  ��  k�  L�  ,�  �  ��  ��  ��  ��  p�  P�  1�  �  ��  ��  ��  ��  s�  S�  3�  �  ��  ��  ��  ��  t�  T�  4�  �  ��  ��  ��  ��  s�  S�  2�  �  ��  ��  ��  ��  p�  P�  /�  �  ��  ��  ��  ��  k�  K�  *�  	�  ��  ��  ��  ��  e�  D�  #�  �  ��  ��  ��  ~�  \�  ;�  �  ��  ؿ  ��  ��  t�  R�  1�  �  �  ̾  ��  ��  h�  F�  $�  �  �  ��  ��  |�  Z�  8�  �  ��  Ҽ  ��  ��  m�  J�  (�  �  �  »  ��  ~�  [�  9�  �  ��  Һ  ��  ��  k�  H�  &�  �  �  ��  ��  y�  V�  4�  �  �  ̸  ��  ��  c�  @�  �  ��  ׷  ��  ��  n�  K�  (�  �  �  ��  ��  x�  U�  2�  �  �  ȵ  ��  ��  ]�  :�  �  �  ϴ  ��  ��  d�  A�  �  ��  ճ  ��  ��  j�  F�  "�  ��  ڲ  ��  ��  n�  J�  &�  �  ޱ  ��  ��  q�  M�  )�  �  �  ��  ��  s�  O�  *�  �  �  ��  ��  s�  O�  *�  �  �  ��  ��  s�  N�  )�  �  ߭  ��  ��  p�  K�  &�  �  ܬ  ��  ��  m�  H�  #�  ��  ث  ��  ��  h�  C�  �  ��  Ӫ  ��  ��  b�  =�  �  �  ̩  ��  ��  [�  5�  �  �  Ĩ  ��  x�  S�  -�  �  �  ��  ��  o�  I�  #�  ��  צ  ��  ��  d�  >�  �  �  ˥  ��  ~�  X�  2�  �  �  ��  ��  q�  K�  $�  ��  ף  ��  ��  c�  <�  �  �  Ȣ  ��  {�  T�  -�  �  ߡ  ��  ��  j�  C�  �  ��  Π  ��  ��  X�  1�  
�  �  ��  ��  m�  E�  �  ��  Ϟ  ��  ��  Y�  1�  
�  �  ��  ��  l�  D�  �  ��  ͜  ��  }�  U�  .�  �  ޛ  ��  ��  f�  >�  �  �  ƚ  ��  v�  N�  &�  ��  ֙  ��  ��  ]�  5�  �  �  ��  ��  k�  C�  �  �  ɗ  ��  x�  P�  '�  ��  ֖  ��  ��  \�  3�  �  �  ��  ��  h�  ?�  �  �  Ĕ  ��  r�  I�   �  ��  Γ  ��  |�  S�  *�  �  ؒ  ��  ��  \�  3�  
�  ��  ��  ��  d�  ;�  �  �  ��  ��  l�  B�  �  �  ŏ  ��  r�  I�  �  ��  ̎  ��  x�  N�  $�  ��  э  ��  }�  S�  )�  ��  Ռ  ��  ��  W�  -�  �  ً  ��  ��  [�  1�  �  ܊  ��  ��  ]�  3�  	�  މ  ��  ��  _�  5�  
�  ��  ��  ��  `�  6�  �  �  ��  ��  a�  6�  �  �  ��  ��  `�  6�  �  ��  ��  ��  _�  4�  	�  ߄  ��  ��  ^�  3�  �  ܃  ��  ��  [�  0�  �  ڂ  ��  ��  X�  -�  �  ց  ��  �  T�  )�  ��  Ҁ  ��  {�  O�  $�  �  �  �  v  J    �~  �~  �~  p~  D~  ~  �}  �}  �}  i}  =}  }  �|  �|  �|  b|  6|  
|  �{  �{  �{  Z{  .{  {  �z  �z  }z  Qz  %z  �y  �y  �y  ty  Hy  y  �x  �x  �x  jx  >x  x  �w  �w  �w  `w  3w  w  �v  �v  �v  Uv  (v  �u  �u  �u  vu  Iu  u  �t  �t  �t  it  =t  t  �s  �s  �s  ]s  0s  s  �r  �r  |r  Or  "r  �q  �q  �q  nq  Aq  q  �p  �p  �p  _p  2p  p  �o  �o  }o  Po  #o  �n  �n  �n  mn  @n  n  �m  �m  �m  ]m  0m  m  �l  �l  zl  Ll  l  �k  �k  �k  hk  :k  k  �j  �j  �j  Vj  (j  �i  �i  �i  qi  Ci  i  �h  �h  �h  ^h  0h  h  �g  �g  xg  Jg  g  �f  �f  �f  df  6f  f  �e  �e  ~e  Pe  !e  �d  �d  �d  id  :d  d  �c  �c  �c  Sc  %c  �b  �b  �b  kb  =b  b  �a  �a  �a  Ta  &a  �`  �`  �`  l`  =`  `  �_  �_  �_  T_  %_  �^  �^  �^  k^  <^  ^  �]  �]  �]  R]  #]  �\  �\  �\  h\  9\  
\  �[  �[  }[  N[  [  �Z  �Z  �Z  cZ  4Z  Z  �Y  �Y  xY  IY  Y  �X  �X  �X  ]X  .X  �W  �W  �W  qW  BW  W  �V  �V  �V  VV  &V  �U  �U  �U  iU  9U  
U  �T  �T  |T  LT  T  �S  �S  �S  _S  /S   S  �R  �R  qR  AR  R  �Q  �Q  �Q  SQ  $Q  �P  �P  �P  eP  5P  P  �O  �O  vO  FO  O  �N  �N  �N  WN  'N  �M  �M  �M  hM  8M  M  �L  �L  xL  HL  L  �K  �K  �K  XK  (K  �J  �J  �J  hJ  8J  J  �I  �I  wI  GI  I  �H  �H  �H  VH  &H  �G  �G  �G  eG  4G  G  �F  �F  sF  CF  F  �E  �E  �E  QE  !E  �D  �D  �D  _D  /D  �C  �C  �C  mC  <C  C  �B  �B  zB  JB  B  �A  �A  �A  WA  &A  �@  �@  �@  d@  3@  @  �?  �?  p?  ??  ?  �>  �>  }>  L>  >  �=  �=  �=  X=  '=  �<  �<  �<  d<  3<  <  �;  �;  o;  ?;  ;  �:  �:  {:  J:  :  �9  �9  �9  U9  $9  �8  �8  �8  `8  /8  �7  �7  �7  k7  :7  	7  �6  �6  u6  D6  6  �5  �5  �5  N5  5  �4  �4  �4  Y4  '4  �3  �3  �3  b3  13   3  �2  �2  l2  ;2  
2  �1  �1  v1  D1  1  �0  �0  0  N0  0  �/  �/  �/  W/  %/  �.  �.  �.  `.  ..  �-  �-  �-  h-  7-  -  �,  �,  q,  ?,  ,  �+  �+  y+  H+  +  �*  �*  �*  P*  *  �)  �)  �)  X)  &)  �(  �(  �(  `(  .(  �'  �'  �'  h'  6'  '  �&  �&  o&  >&  &  �%  �%  w%  E%  %  �$  �$  ~$  L$  $  �#  �#  �#  S#  "#  �"  �"  �"  Z"  )"  �!  �!  �!  a!  0!  �   �   �   h   6      �  �  o  =    �  �  u  C    �  �  |  J    �  �  �  P    �  �  �  V  $  �  �  �  \  *  �  �  �  b  0  �  �  �  h  6    �  �  n  <  
  �  �  t  A    �  �  y  G    �  �    M    �  �  �  R     �  �  �  W  %  �  �  �  ]  *  �  �  �  b  0  �  �  �  g  5    �  �  l  :    �  �  q  ?    �  �  v  D    �  �  {  I    �
  �
  �
  N
  
  �	  �	  �	  S	   	  �  �  �  W  %  �  �  �  \  *  �  �  �  a  /  �  �  �  f  3    �  �  j  8    �  �  o  =    �  �  t  B    �  �  x  F    �   �   }   K      ������������Q������������������U���#���������������Z���(���������������_���,���������������c���1���������������h���6��������������m���;��������������r���?��������������v���D��������������{���I������������������N������������������S���!���������������X���%���������������]���+���������������b���0���������������g���5��������������l���:��������������q���?��������������w���D��������������|���J������������������O������������������U���#���������������Z���(���������������`���.���������������f���4��������������l���:��������������r���@��������������x���F��������������~���L������������������R��� ���������������Y���'���������������_���-���������������f���4��������������m���;���	�����������t���B��������������{���I������������������P������������������X���&���������������_���-���������������g���5��������������n���=��������������v���E��������������~���M������������������U���$���������������^���,���������������f���5��������������o���>��������������x���F������������������P������������������Y���(���������������c���1��� �����������l���;���
�����������v���E������������������O������������������Z���(���������������d���3��������������o���>��������������z���I������������������T���#���������������`���/���������������k���;���
�����������w���F������������������S���"���������������_���.�������Ϳ������l���;������ھ������y���H�����������������U���%�������ļ������c���2������ѻ������q���@������ߺ���������N�����������������\���,�������̸������k���;������ڷ������z���J�����������������Y���)�������ȵ������h���8������ش������x���H�����������������X���(�������Ȳ������h���8���	���ٱ������y���I�����������������Z���*�������˯������k���<������ܮ������}���M�����������������_���0��� ���Ѭ������r���B�����������������U���%�������Ǫ������h���8���	���ک������{���L�����������������_���0������ҧ������t���D�����������������Y���*�������̥������n���?�����������������T���%�������ǣ������i���:������ݢ���������P���"������ġ������g���8���	���۠������}���O��� ������ß������f���7���	���ڞ������}���O��� ������Ý������g���8���
���ۜ���������P���"�������ƛ������i���;������ߚ����������T���&�������ʙ������n���@�����������������Z���,�������З������t���F�����������������a���3������ؕ������|���O���!������Ɣ������j���=�����������������Y���+�������В������v���H�����������������e���8������ݐ����������V���(�������Ώ������t���F�����������������e���8������ލ����������W���*�������Ќ������w���J����������Ë������j���=�����������������^���1������؉���������R���&�������͈������t���G���������������i���=�����������������`���3������ۅ����������V���*�������҄������z���N���"�������ʃ������r���F���������Â������k���?�����������������e���9�����������������_���3���������������Z��.�����~���~���~��U~��*~���}���}���}��}}��R}��&}���|���|���|��z|��O|��$|���{���{���{��w{��L{��!{���z���z���z��vz��Kz�� z���y���y���y��uy��Jy��y���x���x���x��ux��Jx��x���w���w���w��uw��Kw�� w���v���v���v��vv��Lv��"v���u���u���u��xu��Nu��$u���t���t���t��{t��Qt��'t���s���s���s��s��Us��+s��s���r���r���r��Yr��/r��r���q���q���q��^q��5q��q���p���p���p��dp��;p��p���o���o���o��ko��Ao��o���n���n���n��rn��In�� n���m���m���m��{m��Qm��(m���l���l���l���l��[l��2l��	l���k���k���k��ek��<k��k���j���j���j��pj��Gj��j���i���i���i��{i��Si��*i��i���h���h���h��_h��7h��h���g���g���g��mg��Dg��g���f���f���f��{f��Sf��*f��f���e���e���e��be��:e��e���d���d���d��rd��Jd��"d���c���c���c���c��[c��3c��c���b���b���b��mb��Eb��b���a���a���a���a��Xa��1a��	a���`���`���`��l`��E`��`���_���_���_���_��Y_��2_��_���^���^���^��o^��H^��!^���]���]���]���]��_]��8]��]���\���\���\��v\��P\��)\��\���[���[���[��h[��B[��[���Z���Z���Z���Z��[Z��5Z��Z���Y���Y���Y��vY��PY��)Y��Y���X���X���X��kX��EX��X���W���W���W���W��bW��<W��W���V���V���V��V��ZV��4V��V���U���U���U��xU��SU��-U��U���T���T���T��rT��MT��(T��T���S���S���S��nS��IS��$S���R���R���R���R��kR��FR��!R���Q���Q���Q���Q��iQ��DQ��Q���P���P���P���P��hP��CP��P���O���O���O���O��iO��DO�� O���N���N���N���N��jN��FN��"N���M���M���M���M��nM��JM��&M��M���L���L���L��rL��NL��+L��L���K���K���K��xK��TK��1K��K���J���J���J��J��\J��8J��J���I���I���I���I��eI��AI��I���H���H���H���H��oH��LH��)H��H���G���G���G��zG��WG��4G��G���F���F���F���F��dF��BF��F���E���E���E���E��sE��PE��.E��E���D���D���D���D��`D��>D��D���C���C���C���C��qC��PC��.C��C���B���B���B���B��bB��AB��B���A���A���A���A��wA��UA��4A��A���@���@���@���@��k@��J@��(@��@���?���?���?���?��a?��@?��?���>���>���>���>��z>��Y>��8>��>���=���=���=���=��t=��S=��3=��=���<���<���<���<��o<��O<��/<��<���;���;���;���;��m;��M;��-;��;���:���:���:���:��l:��L:��,:��:���9���9���9���9��n9��N9��.9��9���8���8���8���8��q8��Q8��28��8���7���7���7���7��v7��W7��77��7���6���6���6���6��}6��^6��?6�� 6��6���5���5���5���5��g5��H5��*5��5���4���4���4���4��r4��T4��54��4���3���3���3���3��3��a3��C3��%3��3���2���2���2���2��p2��S2��52��2���1���1���1���1���1��d1��F1��)1��1���0���0���0���0��x0��Z0��=0�� 0��0���/���/���/���/��p/��S/��6/��/���.���.���.���.���.��k.��N.��1.��.���-���-���-���-���-��i-��L-��/-��-���,���,���,���,���,��i,��L,��0,��,���+���+���+���+���+��k+��O+��3+��+���*���*���*���*���*��p*��U*��9*��*��*���)���)���)���)��x)��])��B)��&)��)���(���(���(���(���(��h(��M(��2(��(���'���'���'���'���'��u'��Z'��?'��%'��
'���&���&���&���&���&��k&��P&��6&��&��&���%���%���%���%��~%��c%��I%��/%��%���$���$���$���$���$��y$��_$��F$��,$��$���#���#���#���#���#��x#��_#��E#��,#��#���"���"���"���"���"��{"��b"��H"��/"��"���!���!���!���!���!���!��h!��O!��6!��!��!��� ��� ��� ��� ��� ��q ��Y ��@ ��( �� �����������������~��f��N��6���������������������v��^��G��/���� �����������������s��[��D��-����������������������s��\��E��.���������������������x��a��K��4������������������������k��U��>��(����������������������x��b��M��7��!����������������������t��_��J��4����
��������������������v��a��L��7��"����������������������|��g��S��>��*������������������������s��_��K��7��#�������������������������p��]��I��5��"�������������������������t��`��M��:��'������������������������}��j��W��E��2���������������������������z��g��U��C��1���������������������������~��l��Z��I��7��%���������������������������w��f��U��D��3��"���� �����������������������y��i��X��H��7��'������������������������������t��d��S��C��4��$������������������������������w��h��X��I��9��*���������������������������������u��f��W��H��:��+�������
���
���
���
���
���
���
���
���
��~
��o
��a
��S
��E
��7
��)
��
��
���	���	���	���	���	���	���	���	���	���	��v	��h	��[	��M	��@	��2	��%	��	��	��������������������������������{��n��b��U��H��;��/��"����	�����������������������������������v��j��^��R��F��:��.��#������������������������������������������v��k��`��U��I��>��3��(��������������������������������������������~��t��i��_��U��K��@��6��,��"�����������������������������������������������}��t��k��b��X��O��F��=��4��+��"�����������������������������������������������������~��u��m��e��]��U��M��E��=��5��-��%����������������������������������������������������������������z��t��m��f��_��X��Q��K��D��=��7��0��*��#��������	����������������������������������������������������������������������}��w��r��m��g��b��]��X��S��N��I��D��?��:��5��0��+��&��"����������
������� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��} ��z ��w ��t ��q ��n ��k ��i ��f ��c ��` ��^ ��[ ��X ��V ��S ��Q ��N ��L ��I ��G ��E ��B ��@ ��> ��< ��: ��8 ��6 ��4 ��2 ��0 ��. ��, ��* ��( ��' ��% ��# ��" ��  �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��
 ��	 ��	 �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��	 ��	 ��
 �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��  ��" ��# ��% ��' ��( ��* ��, ��. ��0 ��2 ��4 ��6 ��8 ��: ��< ��> ��@ ��B ��E ��G ��I ��L ��N ��Q ��S ��V ��X ��[ ��^ ��` ��c ��f ��i ��k ��n ��q ��t ��w ��z ��} ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ������
����������"��&��+��0��5��:��?��D��I��N��S��X��]��b��g��m��r��w��}����������������������������������������������������������������������	��������#��*��0��7��=��D��K��Q��X��_��f��m��t��z����������������������������������������������������������������%��-��5��=��E��M��U��]��e��m��u��~�����������������������������������������������������"��+��4��=��F��O��X��b��k��t��}�����������������������������������������������"��,��6��@��K��U��_��i��t��~��������������������������������������������(��3��>��I��U��`��k��v������������������������������������������#��.��:��F��R��^��j��v�����������������������������������	����"��/��;��H��U��b��n��{��������������������������������	��	��%	��2	��@	��M	��[	��h	��v	���	���	���	���	���	���	���	���	���	���	��
��
��)
��7
��E
��S
��a
��o
��~
���
���
���
���
���
���
���
���
���
������+��:��H��W��f��u���������������������������������*��9��I��X��h��w������������������������������$��4��C��S��d��t������������������������������'��7��H��X��i��y����������������������� ����"��3��D��U��f��w���������������������������%��7��I��Z��l��~���������������������������1��C��U��g��z���������������������������2��E��W��j��}������������������������'��:��M��`��t�������������������������"��5��I��]��p�������������������������#��7��K��_��s������������������������*��>��S��g��|����������������������"��7��L��a��v��������������������
����4��J��_��t����������������������!��7��M��b��x����������������������(��>��U��k������������������������4��K��a��x���������������������.��E��\��s����������������������-��D��[��s����������������� ����/��G��^��v���������������������6��N��f��~����������������� ��( ��@ ��Y ��q ��� ��� ��� ��� ��� ��!��!��6!��O!��h!���!���!���!���!���!���!��"��/"��H"��b"��{"���"���"���"���"���"��#��,#��E#��_#��x#���#���#���#���#���#��$��,$��F$��_$��y$���$���$���$���$���$��%��/%��I%��c%��~%���%���%���%���%��&��&��6&��P&��k&���&���&���&���&���&��
'��%'��?'��Z'��u'���'���'���'���'���'��(��2(��M(��h(���(���(���(���(���(��)��&)��B)��])��x)���)���)���)���)��*��*��9*��U*��p*���*���*���*���*���*��+��3+��O+��k+���+���+���+���+���+��,��0,��L,��i,���,���,���,���,���,��-��/-��L-��i-���-���-���-���-���-��.��1.��N.��k.���.���.���.���.���.��/��6/��S/��p/���/���/���/���/��0�� 0��=0��Z0��x0���0���0���0���0��1��)1��F1��d1���1���1���1���1���1��2��52��S2��p2���2���2���2���2��3��%3��C3��a3��3���3���3���3���3��4��54��T4��r4���4���4���4���4��5��*5��H5��g5���5���5���5���5��6�� 6��?6��^6��}6���6���6���6���6��7��77��W7��v7���7���7���7���7��8��28��Q8��q8���8���8���8���8��9��.9��N9��n9���9���9���9���9��:��,:��L:��l:���:���:���:���:��;��-;��M;��m;���;���;���;���;��<��/<��O<��o<���<���<���<���<��=��3=��S=��t=���=���=���=���=��>��8>��Y>��z>���>���>���>���>��?��@?��a?���?���?���?���?��@��(@��J@��k@���@���@���@���@��A��4A��UA��wA���A���A���A���A��B��AB��bB���B���B���B���B��C��.C��OC��qC���C���C���C���C��D��>D��`D���D���D���D���D��E��.E��PE��sE���E���E���E���E��F��BF��dF���F���F���F���F��G��5G��WG��zG���G���G���G��H��)H��LH��oH���H���H���H���H��I��AI��eI���I���I���I���I��J��8J��\J��J���J���J���J��K��1K��UK��xK���K���K���K��L��+L��NL��rL���L���L���L��M��&M��JM��nM���M���M���M���M��"N��FN��jN���N���N���N���N�� O��DO��iO���O���O���O���O��P��CP��hP���P���P���P���P��Q��DQ��iQ���Q���Q���Q���Q��!R��FR��kR���R���R���R���R��$S��IS��nS���S���S���S��T��(T��MT��rT���T���T���T��U��-U��SU��xU���U���U���U��V��4V��ZV��V���V���V���V��W��<W��bW���W���W���W���W��X��EX��kX���X���X���X��Y��)Y��PY��vY���Y���Y���Y��Z��5Z��[Z���Z���Z���Z���Z��[��B[��h[���[���[���[��\��)\��P\��v\���\���\���\��]��8]��_]���]���]���]���]��!^��H^��o^���^���^���^��_��2_��Y_���_���_���_���_��`��E`��l`���`���`���`��	a��1a��Xa���a���a���a���a��b��Eb��mb���b���b���b��c��3c��[c���c���c���c���c��"d��Jd��rd���d���d���d��e��:e��be���e���e���e��f��*f��Sf��{f���f���f���f��g��Dg��mg���g���g���g��h��7h��_h���h���h���h��i��*i��Si��{i���i���i���i��j��Gj��pj���j���j���j��k��<k��ek���k���k���k��	l��2l��[l���l���l���l���l��(m��Rm��{m���m���m���m�� n��In��rn���n���n���n��o��Ao��ko���o���o���o��p��;p��dp���p���p���p��q��4q��^q���q���q���q��r��/r��Yr���r���r���r��s��+s��Us��s���s���s���s��'t��Qt��{t���t���t���t��$u��Nu��xu���u���u���u��"v��Lv��vv���v���v���v�� w��Kw��uw���w���w���w��x��Jx��ux���x���x���x��y��Jy��uy���y���y���y�� z��Kz��vz���z���z���z��!{��L{��w{���{���{���{��$|��O|��z|���|���|���|��&}��R}��}}���}���}���}��*~��U~���~���~���~����.��Z��������������3���_�����������������9���e�����������������?���k�������Â��������F���r�������ʃ������"���N���z�������҄������*���V�����������ۅ�����3���`�����������������=���i���������������G���t�������͈������&���R����������؉�����1���^�����������������=���j�������Ë���������J���w�������Ќ������*���W�����������ލ�����8���e�����������������F���t�������Ώ������(���V�����������ݐ�����8���e�����������������H���v�������В������+���Y�����������������=���j�������Ɣ�����!���O���|�������ؕ�����3���a�����������������F���t�������З������,���Z�����������������@���n�������ʙ������&���T�����������ߚ�����;���i�������ƛ������"���P����������ۜ��
���8���g�������Ý����� ���O���}�������ڞ��	���7���f�������ß����� ���O���}�������۠��	���8���g�������ġ�����"���P����������ݢ�����:���i�������ǣ������%���T�����������������?���n�������̥������*���Y�����������������D���t�������ҧ�����0���`�����������������L���{�������ک��	���8���h�������Ǫ������%���U�����������������B���r�������Ѭ�� ���0���_�����������������M���}�������ܮ�����<���k�������˯������*���Z�����������������I���y�������ٱ��	���8���h�������Ȳ������(���X�����������������H���x�������ش�����8���h�������ȵ������)���Y�����������������J���z�������ڷ�����;���k�������̸������,���\�����������������N����������ߺ�����@���q�������ѻ�����2���c�������ļ������%���U�����������������H���y�������ھ�����;���l�������Ϳ������.���_���������������"���S������������������F���w�����������
���;���k���������������/���`���������������#���T������������������I���z��������������>���o��������������3���d���������������(���Z������������������O������������������E���v�����������
���;���l����������� ���1���c���������������(���Y������������������P������������������G���x��������������>���o��������������5���f���������������,���^���������������$���U������������������M���~��������������E���v��������������=���n��������������5���g���������������-���_���������������&���X������������������P������������������I���{��������������B���t�����������	���;���m��������������4���f���������������-���_���������������'���Y��������������� ���R������������������L���~��������������F���x��������������@���r��������������:���l��������������4���f���������������.���`���������������(���Z���������������#���U������������������O������������������J���|��������������D���w��������������?���q��������������:���l��������������5���g���������������0���b���������������+���]���������������%���X���������������!���S������������������N������������������I���{��������������D���v��������������?���r��������������;���m��������������6���h���������������1���c���������������,���_���������������(���Z���������������#���U������������������Q���������������   K   }   �   �     F  x  �  �    B  t  �  �    =  o  �  �    8  j  �  �    3  f  �  �  �  /  a  �  �  �  *  \  �  �  �  %  W  �  �  �   	  S	  �	  �	  �	  
  N
  �
  �
  �
    I  {  �  �    D  v  �  �    ?  q  �  �    :  l  �  �    5  g  �  �  �  0  b  �  �  �  *  ]  �  �  �  %  W  �  �  �     R  �  �  �    M    �  �    G  y  �  �    A  s  �  �  
  <  n  �  �    6  h  �  �  �  0  b  �  �  �  *  \  �  �  �  $  V  �  �  �    P  �  �  �    J  |  �  �    C  u  �  �    =  o  �  �     6   h   �   �   �   0!  a!  �!  �!  �!  )"  Z"  �"  �"  �"  "#  S#  �#  �#  �#  $  L$  ~$  �$  �$  %  E%  w%  �%  �%  &  >&  o&  �&  �&  '  6'  h'  �'  �'  �'  .(  `(  �(  �(  �(  &)  X)  �)  �)  �)  *  P*  �*  �*  �*  +  H+  y+  �+  �+  ,  ?,  q,  �,  �,  -  7-  h-  �-  �-  �-  ..  `.  �.  �.  �.  %/  W/  �/  �/  �/  0  N0  0  �0  �0  1  D1  v1  �1  �1  
2  ;2  l2  �2  �2   3  13  b3  �3  �3  �3  '4  Y4  �4  �4  �4  5  O5  �5  �5  �5  6  D6  u6  �6  �6  	7  :7  k7  �7  �7  �7  /8  `8  �8  �8  �8  $9  U9  �9  �9  �9  :  J:  {:  �:  �:  ;  ?;  o;  �;  �;  <  3<  d<  �<  �<  �<  '=  X=  �=  �=  �=  >  L>  }>  �>  �>  ?  ??  p?  �?  �?  @  3@  d@  �@  �@  �@  &A  WA  �A  �A  �A  B  JB  zB  �B  �B  C  <C  mC  �C  �C  �C  /D  _D  �D  �D  �D  !E  QE  �E  �E  �E  F  CF  sF  �F  �F  G  4G  eG  �G  �G  �G  &H  VH  �H  �H  �H  I  GI  wI  �I  �I  J  8J  hJ  �J  �J  �J  (K  XK  �K  �K  �K  L  HL  xL  �L  �L  M  8M  hM  �M  �M  �M  'N  WN  �N  �N  �N  O  FO  vO  �O  �O  P  5P  eP  �P  �P  �P  $Q  SQ  �Q  �Q  �Q  R  AR  qR  �R  �R   S  /S  _S  �S  �S  �S  T  LT  |T  �T  �T  
U  9U  iU  �U  �U  �U  &V  VV  �V  �V  �V  W  BW  qW  �W  �W  �W  .X  ]X  �X  �X  �X  Y  IY  xY  �Y  �Y  Z  4Z  cZ  �Z  �Z  �Z  [  N[  }[  �[  �[  
\  9\  h\  �\  �\  �\  #]  R]  �]  �]  �]  ^  <^  k^  �^  �^  �^  %_  T_  �_  �_  �_  `  =`  l`  �`  �`  �`  &a  Ta  �a  �a  �a  b  =b  kb  �b  �b  �b  %c  Sc  �c  �c  �c  d  :d  id  �d  �d  �d  !e  Pe  ~e  �e  �e  f  6f  df  �f  �f  �f  g  Jg  xg  �g  �g  h  0h  ^h  �h  �h  �h  i  Ci  qi  �i  �i  �i  (j  Vj  �j  �j  �j  k  :k  hk  �k  �k  �k  l  Ll  zl  �l  �l  m  0m  ]m  �m  �m  �m  n  @n  mn  �n  �n  �n  #o  Po  }o  �o  �o  p  2p  _p  �p  �p  �p  q  Aq  nq  �q  �q  �q  "r  Or  |r  �r  �r  s  0s  ]s  �s  �s  �s  t  =t  it  �t  �t  �t  u  Iu  vu  �u  �u  �u  (v  Uv  �v  �v  �v  w  4w  `w  �w  �w  �w  x  >x  jx  �x  �x  �x  y  Hy  ty  �y  �y  �y  %z  Qz  }z  �z  �z  {  .{  Z{  �{  �{  �{  
|  6|  b|  �|  �|  �|  }  =}  i}  �}  �}  �}  ~  D~  p~  �~  �~  �~    J  v  �  �  �  $�  O�  {�  ��  Ҁ  ��  )�  T�  �  ��  ց  �  -�  X�  ��  ��  ڂ  �  0�  [�  ��  ��  ܃  �  3�  ^�  ��  ��  ߄  	�  4�  _�  ��  ��  ��  �  6�  `�  ��  ��  �  �  6�  a�  ��  ��  �  �  6�  `�  ��  ��  ��  
�  5�  _�  ��  ��  މ  	�  3�  ]�  ��  ��  ܊  �  1�  [�  ��  ��  ً  �  -�  W�  ��  ��  Ռ  ��  )�  S�  }�  ��  э  ��  $�  N�  x�  ��  ̎  ��  �  I�  r�  ��  ŏ  �  �  B�  l�  ��  ��  �  �  ;�  d�  ��  ��  ��  
�  3�  \�  ��  ��  ؒ  �  *�  S�  |�  ��  Γ  ��   �  I�  r�  ��  Ĕ  �  �  ?�  h�  ��  ��  �  �  3�  \�  ��  ��  ֖  ��  '�  P�  x�  ��  ɗ  �  �  C�  k�  ��  ��  �  �  5�  ]�  ��  ��  ֙  ��  &�  N�  v�  ��  ƚ  �  �  >�  f�  ��  ��  ޛ  �  .�  U�  }�  ��  ͜  ��  �  D�  k�  ��  ��  �  
�  1�  Y�  ��  ��  Ϟ  ��  �  E�  m�  ��  ��  �  
�  1�  X�  �  ��  Π  ��  �  C�  j�  ��  ��  ߡ  �  -�  T�  {�  ��  Ȣ  �  �  <�  c�  ��  ��  ף  ��  $�  K�  q�  ��  ��  �  �  2�  X�  ~�  ��  ˥  �  �  >�  d�  ��  ��  צ  ��  #�  I�  o�  ��  ��  �  �  -�  S�  x�  ��  Ĩ  �  �  5�  [�  ��  ��  ̩  �  �  =�  b�  ��  ��  Ӫ  ��  �  C�  h�  ��  ��  ث  ��  #�  H�  m�  ��  ��  ܬ  �  &�  K�  p�  ��  ��  ߭  �  )�  N�  s�  ��  ��  �  �  *�  O�  s�  ��  ��  �  �  *�  O�  s�  ��  ��  �  �  )�  M�  q�  ��  ��  ޱ  �  &�  J�  n�  ��  ��  ڲ  ��  "�  F�  j�  ��  ��  ճ  ��  �  A�  d�  ��  ��  ϴ  �  �  :�  ]�  ��  ��  ȵ  �  �  2�  U�  x�  ��  ��  �  �  (�  K�  n�  ��  ��  ׷  ��  �  @�  c�  ��  ��  ̸  �  �  4�  V�  y�  ��  ��  �  �  &�  H�  k�  ��  ��  Һ  ��  �  9�  [�  ~�  ��  »  �  �  (�  J�  m�  ��  ��  Ҽ  ��  �  8�  Z�  |�  ��  ��  �  �  $�  F�  h�  ��  ��  ̾  �  �  1�  R�  t�  ��  ��  ؿ  ��  �  ;�  \�  ~�  ��  ��  ��  �  #�  D�  e�  ��  ��  ��  ��  	�  *�  K�  k�  ��  ��  ��  ��  �  /�  P�  p�  ��  ��  ��  ��  �  2�  S�  s�  ��  ��  ��  ��  �  4�  T�  t�  ��  ��  ��  ��  �  3�  S�  s�  ��  ��  ��  ��  �  1�  P�  p�  ��  ��  ��  ��  �  ,�  L�  k�  ��  ��  ��  ��  �  &�  E�  d�  ��  ��  ��  ��  ��  �  =�  [�  z�  ��  ��  ��  ��  �  2�  Q�  o�  ��  ��  ��  ��  �  &�  D�  b�  ��  ��  ��  ��  ��  �  6�  T�  r�  ��  ��  ��  ��  �  %�  C�  `�  ~�  ��  ��  ��  ��  �  0�  M�  k�  ��  ��  ��  ��  ��  �  8�  V�  s�  ��  ��  ��  ��  �  !�  >�  [�  x�  ��  ��  ��  ��  �  %�  B�  ^�  {�  ��  ��  ��  ��  
�  &�  B�  _�  {�  ��  ��  ��  ��  �  %�  A�  ]�  y�  ��  ��  ��  ��  �   �  <�  X�  t�  ��  ��  ��  ��  ��  �  5�  Q�  l�  ��  ��  ��  ��  ��  �  ,�  G�  b�  }�  ��  ��  ��  ��  �  �  :�  U�  p�  ��  ��  ��  ��  ��  �  +�  F�  `�  {�  ��  ��  ��  ��  ��  �  4�  N�  h�  ��  ��  ��  ��  ��  �  �  9�  S�  m�  ��  ��  ��  ��  ��  �  !�  ;�  T�  n�  ��  ��  ��  ��  ��  �   �  9�  S�  l�  ��  ��  ��  ��  ��  �  �  5�  N�  g�  �  ��  ��  ��  ��  ��  �  -�  E�  ^�  v�  ��  ��  ��  ��  ��  	�  !�  :�  R�  j�  ��  ��  ��  ��  ��  ��  �  *�  B�  Z�  r�  ��  ��  ��  ��  ��   �  �  /�  G�  ^�  v�  ��  ��  ��  ��  ��  �  �  0�  G�  _�  v�  ��  ��  ��  ��  ��  ��  �  -�  D�  [�  q�  ��  ��  ��  ��  ��  ��  �  &�  <�  R�  i�  �  ��  ��  ��  ��  ��  �  �  0�  F�  \�  r�  ��  ��  ��  ��  ��  ��  
�   �  6�  K�  a�  v�  ��  ��  ��  ��  ��  ��  �  !�  6�  K�  `�  u�  ��  ��  ��  ��  ��  ��  �  �  1�  F�  [�  o�  ��  ��  ��  ��  ��  ��  ��  �  (�  <�  P�  d�  y�  ��  ��  ��  ��  ��  ��  �  �  -�  A�  T�  h�  |�  ��  ��  ��  ��  ��  ��  �  �  ,�  ?�  S�  f�  y�  ��  ��  ��  ��  ��  ��  ��  �  %�  8�  K�  ^�  q�  ��  ��  ��  ��  ��  ��  ��  �  �  +�  =�  O�  b�  t�  ��  ��  ��  ��  ��  ��  ��  �  �  )�  ;�  M�  _�  q�  ��  ��  ��  ��  ��  ��  ��  ��  �  !�  2�  C�  U�  f�  w�  ��  ��  ��  ��  ��  ��  ��   �  �  "�  3�  D�  T�  e�  v�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  +�  <�  L�  \�  l�  |�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  +�  ;�  K�  Z�  j�  y�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  "�  1�  @�  O�  ^�  m�  |�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  ,�  ;�  I�  X�  f�  t�  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  +�  8�  F�  T�  b�  o�  }�  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  *�  7�  D�  Q�  ^�  k�  x�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  (�  5�  A�  M�  Z�  f�  r�  ~�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  #�  /�  ;�  F�  Q�  ]�  h�  s�  �  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  #�  .�  9�  C�  N�  X�  c�  m�  x�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  #�  -�  6�  @�  J�  S�  ]�  f�  p�  y�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  �  %�  .�  6�  ?�  H�  P�  X�  a�  i�  r�  z�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  	�  �  �   �  (�  /�  6�  >�  E�  L�  T�  [�  b�  i�  p�  w�  �  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  	�  �  �  �  "�  (�  .�  4�  :�  @�  F�  K�  Q�  W�  ]�  b�  h�  m�  s�  x�  ~�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  �  �  �  �  �  !�  %�  )�  -�  1�  5�  9�  =�  A�  E�  H�  L�  P�  S�  W�  [�  ^�  b�  e�  i�  l�  o�  s�  v�  y�  |�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ����Ś��x��|{���C�����j7�U)R��f���v��ԃ��������l��)��P��u���r���y����$���g��!]��*��z���C����������������B�������B��"���;�������7��NH���I���=��!%��� ��a������UU���	��n���W[��*���Q���D!��\����1��Z����-��Ĥ��N������9���W��R���G��w�������'���{��v������9i����������B��C�����������G�������������W2��Di��ў��	�������7��3h�������������2��]J���t��ם��6�������_��6:��C_����������������x��A.��fN���m��ڌ��1�������/���������:���U���p������u���ý�������������� 6���L��Zc��{y��A�������ƹ��������������
��l���1���D��<W���i���{������+�����������u������w���������K#���2��B��5Q��`���n��S}������ə����������"����������������������K�����*��F6��OB��3N���Y���e��q��e|������������������:���Խ��O��������������������������,���!��+��g4���=���F���O���X���a��Lj���r���{��	���r���Ɣ�����/���E���H���6��������������0�������>����������N���������������$���+��~2��E9���?���F��@M���S��GZ���`��g��hm���s���y�����(���7���9���/����������ĩ������@����������!�������)����������a�����������8���k�������� ������
��������������w#��H(��-���1���6��4;���?��vD��	I���M��R���V��[��p_���c��-h���l���p��u��Jy��~}������х��������������!����������������ŭ������q���>����������~���2�����������(�������Z�������s�������w�������c�������:�����������T ��������>
�����������0��`������ ���#���&��*��-��+0��53��;6��<9��9<��2?��&B��E��H���J���M���P���S��\V��.Y���[���^���a��Qd��g���i���l��4o���q���t��8w���y��}|��������I���ۆ��j�������~�������������|������g���ן��E����������z���۫��8����������?�������߹��+���s�����������<���y����������� ���Q�������������������#���D���d����������������������������������
������������������
��� ���������������	��������n��R��3�������������z��O��" ���!���#���%��X'�� )���*���,��n.��.0���1���3��e5��7���8���:��><���=���?��MA���B���D��LF���G���I��;K���L��|N��P���Q��QS���T���V��X���Y��=[���\��]^���_��wa��c���d��f���g��i���j��l���m��o���p��r���s��u��{v���w��dy���z��G|���}��$����������f���΄��5�����������b���ċ��$����������=����������K�����������M����������C����������/���{���ƣ�����X����������+���n����������3���r����������)���d�������ַ�����D���y�������������D���t���������������)���T���~������������������@���c����������������������&���C���_���z�����������������������
������3���F���X���i���y�������������������������������������������������������������
������������������
���������  ��� ���������������������������	���
��������u��e��U��D��3�� ����������������������u��\��C��)�������������� ���!��b"��C#��#$��%���%���&���'��{(��W)��3*��+���+���,���-��u.��M/��%0���0���1���2��}3��R4��&5���5���6���7��q8��B9��:���:���;���<��O=��>���>���?���@��NA��B���B���C��wD��@E��	F���F���G��^H��%I���I���J��tK��8L���L���M���N��DO��P���P���Q��HR��S���S���T��CU��V���V��{W��7X���X���Y��iZ��#[���[���\��P]��^���^��x_��/`���`���a��Rb��c���c��pd��$e���e���f��=g���g���h��Si��j���j��dk��l���l��rm�� n���n��{o��(p���p���q��-r���r���s��.t���t���u��,v���v��~w��&x���x��uy��z���z��i{��|���|��Z}���}���~��G���������0���Ӂ��u����������Y�����������:���ن��y����������T����������,���ɋ��e����������8���ӎ��n����������<���Ց��n����������7���Δ��f�����������)�������U����������������<���Л��d������������������@���ҟ��c������������������4���ģ��S������p������������������5�������N���ک��f������}�����������������1�������D���ί��V���߰��g������w�������������������������%�������0�������:�������C���ǹ��K���κ��R���ջ��W���ڼ��\���޽��`������b������d�������e�������e�������c�������a�������^�������Z�������U�������O�������H�������@�������8�������.�������#�������������������������w�������i�������Y�������I�������8�������&������������������u�������`�������J�������3�����������������w�������^�������D�������(����������~�������a�������C�������%����������u�������U�������4������������������]�������9������������������\�������6����������{�������S�������*������� ���k�������@�����������������S�������&�����������a�������2����������k�������:�������	���p�������>����������r�������>�������
���p�������;����������j�������3 ��� ��� ��_�����'��������Q�������{�����@�������g�����*��������O�����	��r	���	��4
���
���
��U�������u�����4��������R�������o�����,��������F�������_�������x�����2��������H�������]�������q�����(��������:��������K����� ��Z�������i�������v�����)��������5��������? ��� ��� ��I!���!���!��Q"���"��#��Y#���#��$��_$���$��%��d%���%��&��h&���&��'��l'���'��(��n(���(��)��o)���)��*��o*���*��+��o+���+��,��m,���,��-��j-���-��.��g.���.��/��b/���/��	0��\0���0��1��V1���1���1��O2���2���2��F3���3���3��=4���4���4��35���5���5��(6��y6���6��7��m7���7��8��`8���8��9��R9���9���9��C:���:���:��4;���;���;��#<��s<���<��=��a=���=�� >��O>���>���>��;?���?���?��'@��v@���@��A��aA���A���A��KB���B���B��4C���C���C��D��jD���D��E��QE���E���E��8F���F���F��G��jG���G��H��OH���H���H��3I��I���I��J��bJ���J���J��DK���K���K��&L��qL���L��M��QM���M���M��1N��|N���N��O��[O���O���O��9P���P���P��Q��`Q���Q���Q��=R���R���R��S��bS���S���S��=T���T���T��U��`U���U���U��9V���V���V��W��ZW���W���W��2X��zX���X��	Y��QY���Y���Y��'Z��oZ���Z���Z��D[���[���[��\��`\���\���\��4]��{]���]��^��N^���^���^�� _��g_���_���_��8`��~`���`��
a��Oa���a���a�� b��eb���b���b��5c��zc���c��d��Id���d���d��e��\e���e���e��)f��nf���f���f��:g��~g���g��h��Kh���h���h��i��Zi���i���i��$j��hj���j���j��2k��uk���k���k��>l���l���l��m��Jm���m���m��n��Un���n���n��o��^o���o���o��%p��gp���p���p��-q��oq���q���q��4r��vr���r���r��;s��|s���s���s��@t���t���t��u��Eu���u���u��v��Hv���v���v��
w��Kw���w���w��x��Mx���x���x��y��Ny���y���y��z��Oz���z���z��{��N{���{���{��|��M|���|���|��}��K}���}���}��~��H~���~���~����D�����������?���~�����������:���y�����������4���s����������-���l����������&���d��������������\�������ׅ�����R�������Ά�����H�������Ç�����>���{�����������3���p����������'���d�������݊�����W�������Ћ�����I�������������;���w�����������,���h�������������Y�������я�����H���������������7���s����������&���a�������ؒ�����O�������œ�����<���w����������(���c�������ٕ�����O�������Ė������:���u����������$���_�������Ԙ�����I���������������2���l��������������T�������ț�����<���v����������$���]�������ѝ��
���D���~����������*���d�������֟�����I���������������.���g�������١�����K���������������/���h�������٣�����K���������������.���f�������ץ�����H��������������*���b�������ӧ�����C���{����������#���[�������˩�����;���s�������������R�������«������1���i�������ج�����G�������������%���\�������ˮ�����:���q�������߯�����N��������������*���a�������ϱ�����=���t�������������O��������������*���a�������δ�����;���r�������ߵ�����L��������������%���[�������ȷ������4���k�������׸�����C���y�������������R��������������)���_�������˻�����7���l�������ؼ�����C���y�������������O��������������%���[�������ƿ������1���f��������������;���q��������������F���{��������������O���������������#���X���������������,���a����������� ���5���i��������������=���q��������������D���y��������������K������������������R���������������#���X���������������)���^���������������/���c����������� ���4���h��������������8���l�����������	���=���q��������������A���t��������������D���x��������������G���{��������������J���~��������������M������������������O������������������Q������������������R��������������� ���S���������������!���T���������������"���U���������������"���U���������������"���U���������������"���U���������������"���U���������������!���T��������������� ���S������������������R������������������P������������������O������������������M������������������K���~��������������I���{��������������F���y��������������D���v��������������A���s��������������>���p��������������;���m��������������8���j��������������4���g���������������1���c���������������-���_���������������)���\���������������%���X���������������!���T������������������P������������������K���~��������������G���y��������������C���u��������������>���q��������������:���l��������������5���h���������������1���c���������������,���_���������������(���Z���������������#���U������������������Q���������������   K   }   �   �     F  x  �  �    B  t  �  �    =  o  �  �    8  k  �  �    4  f  �  �  �  /  a  �  �  �  +  ]  �  �  �  &  Y  �  �  �  "	  T	  �	  �	  �	  
  P
  �
  �
  �
    L  ~  �  �    H  z  �  �    C  v  �  �    @  r  �  �  	  <  n  �  �    8  j  �  �    4  g  �  �  �  1  c  �  �  �  .  `  �  �  �  *  ]  �  �  �  '  Z  �  �  �  $  W  �  �  �  "  T  �  �  �    R  �  �  �    P  �  �  �    M  �  �  �    L  ~  �  �    J  }  �  �    H  {  �  �    G  z  �  �    F  y  �  �     E   x   �   �   !  E!  x!  �!  �!  "  D"  x"  �"  �"  #  D#  x#  �#  �#  $  E$  x$  �$  �$  %  E%  x%  �%  �%  &  F&  y&  �&  �&  '  G'  z'  �'  �'  (  H(  |(  �(  �(  )  J)  ~)  �)  �)  *  L*  �*  �*  �*  +  N+  �+  �+  �+  ,  Q,  �,  �,  �,   -  T-  �-  �-  �-  $.  X.  �.  �.  �.  '/  [/  �/  �/  �/  +0  _0  �0  �0  �0  01  d1  �1  �1   2  52  i2  �2  �2  3  :3  n3  �3  �3  4  ?4  t4  �4  �4  5  E5  z5  �5  �5  6  L6  �6  �6  �6  7  S7  �7  �7  �7  %8  Z8  �8  �8  �8  -9  b9  �9  �9   :  5:  j:  �:  �:  	;  >;  s;  �;  �;  <  G<  |<  �<  �<  =  P=  �=  �=  �=  %>  Z>  �>  �>  �>  /?  e?  �?  �?  @  :@  p@  �@  �@  A  FA  {A  �A  �A  B  QB  �B  �B  �B  (C  ^C  �C  �C  �C  5D  kD  �D  �D  E  CE  xE  �E  �E  F  QF  �F  �F  �F  )G  _G  �G  �G  H  8H  nH  �H  �H  I  HI  ~I  �I  �I  !J  XJ  �J  �J  �J  2K  iK  �K  �K  L  CL  zL  �L  �L  M  UM  �M  �M  �M  1N  hN  �N  �N  O  DO  {O  �O  �O  !P  XP  �P  �P  �P  5Q  lQ  �Q  �Q  R  JR  �R  �R  �R  (S  _S  �S  �S  T  >T  vT  �T  �T  U  UU  �U  �U  �U  5V  mV  �V  �V  W  MW  �W  �W  �W  -X  fX  �X  �X  Y  GY  Y  �Y  �Y  )Z  aZ  �Z  �Z  [  D[  |[  �[  �[  '\  _\  �\  �\  
]  C]  |]  �]  �]  '^  `^  �^  �^  _  E_  ~_  �_  �_  *`  c`  �`  �`  a  Ia  �a  �a  �a  /b  ib  �b  �b  c  Pc  �c  �c  �c  8d  rd  �d  �d   e  Ze  �e  �e  f  Cf  }f  �f  �f  ,g  gg  �g  �g  h  Qh  �h  �h  i  <i  vi  �i  �i  'j  bj  �j  �j  k  Nk  �k  �k  �k  ;l  vl  �l  �l  (m  cm  �m  �m  n  Qn  �n  �n  o  @o  |o  �o  �o  /p  kp  �p  �p  q  \q  �q  �q  r  Lr  �r  �r  s  >s  zs  �s  �s  0t  mt  �t  �t  #u  `u  �u  �u  v  Sv  �v  �v  
w  Hw  �w  �w  �w  =x  zx  �x  �x  2y  py  �y  �y  )z  gz  �z  �z   {  ^{  �{  �{  |  V|  �|  �|  }  O}  �}  �}  
~  I~  �~  �~    C  �  �  �  >�  }�  ��  ��  :�  y�  ��  ��  7�  v�  ��  ��  4�  t�  ��  �  3�  r�  ��  �  2�  r�  ��  �  2�  r�  ��  �  2�  s�  ��  �  4�  t�  ��  ��  6�  w�  ��  ��  9�  z�  ��  ��  >�  �  ��  �  C�  ��  Ō  �  H�  ��  ̍  �  O�  ��  ӎ  �  W�  ��  ۏ  �  _�  ��  �  &�  i�  ��  �  1�  s�  ��  ��  <�  �    �  H�  ��  Δ  �  U�  ��  ܕ  �  c�  ��  �  .�  r�  ��  ��  =�  ��  Ƙ  
�  N�  ��  י  �  `�  ��  �  .�  r�  ��  ��  A�  ��  ˜  �  V�  ��  ��  &�  k�  ��  ��  <�  ��  ȟ  �  S�  ��  �  &�  l�  ��  ��  ?�  ��  ̢  �  Y�  ��  �  .�  u�  ��  �  J�  ��  ٥   �  h�  ��  ��  >�  ��  Χ  �  ^�  ��  �  6�  ~�  ǩ  �  X�  ��  �  2�  z�  ë  �  U�  ��  �  1�  z�  í  �  V�  ��  �  3�  }�  ǯ  �  [�  ��  �  :�  ��  ϱ  �  d�  ��  ��  D�  ��  ڳ  &�  q�  ��  �  S�  ��  �  6�  ��  Ͷ  �  e�  ��  ��  J�  ��  �  /�  |�  ȹ  �  b�  ��  ��  I�  ��  �  1�  �  ̼  �  h�  ��  �  Q�  ��  �  <�  ��  ٿ  '�  v�  ��  �  b�  ��   �  P�  ��  ��  >�  ��  ��  -�  |�  ��  �  l�  ��  �  ]�  ��  ��  O�  ��  ��  B�  ��  ��  5�  ��  ��  *�  {�  ��  �  q�  ��  �  g�  ��  �  _�  ��  �  W�  ��  ��  P�  ��  ��  J�  ��  ��  F�  ��  ��  B�  ��  ��  ?�  ��  ��  =�  ��  ��  ;�  ��  ��  ;�  ��  ��  <�  ��  ��  >�  ��  ��  A�  ��  ��  E�  ��  ��  J�  ��  ��  P�  ��  ��  W�  ��  �  _�  ��  �  h�  ��  �  r�  ��  $�  }�  ��  0�  ��  ��  =�  ��  ��  K�  ��   �  [�  ��  �  k�  ��  !�  }�  ��  4�  ��  ��  G�  ��  ��  \�  ��  �  q�  ��  +�  ��  ��  C�  ��  ��  \�  ��  �  v�  ��  3�  ��  ��  O�  ��  �  l�  ��  +�  ��  ��  K�  ��  �  l�  ��  -�  ��  ��  P�  ��  �  t�  ��  7�  ��  ��  ^�  ��  #�  ��  ��  K�  ��  �  u�  ��  =�  ��  �  i�  ��  2  �  �  ` � + � � \ � ( � � [ � ) � � ^ � - � � f	 �	 7
 �
  q � D �  � � U � * �   k � B �  � � ^ � 7 �  ~ � Y � 5 �  � � ] � < �  � � k � L � . �  � � e  �  J! �! /" �" # �# �# p$ �$ X% �% A& �& +' �' ( �( ) w) �) d* �* Q+ �+ @, �, /- �- . �. / �/ 0 {0 �0 n1 �1 b2 �2 W3 �3 M4 �4 D5 �5 <6 �6 47 �7 .8 �8 (9 �9 $: �:  ; �; < �< = �= > �> ? �? @ �@ A �A "B �B &C �C +D �D 2E �E 9F �F AG �G KH �H UI �I `J �J mK �K zL M �M N �N !O �O 2P �P EQ �Q XR �R mS �S �T U �U &V �V ?W �W XX �X sY Z �Z [ �[ <\ �\ [] �] |^ _ �_ .` �` Ra �a vb 	c �c 0d �d Xe �e �f g �g Ah �h mi j �j 2k �k al �l �m +n �n ^o �o �p -q �q cr �r �s 7t �t qu v �v Jw �w �x 'y �y fz { �{ H| �| �} -~ �~ s � �� ]� � �� L� � �� =� � �� 2� ڇ �� +� ԉ ~� '� ҋ |� '� Ӎ � +� ؏ �� 2� �� �� =� � �� L� �� �� _� � Ø u� (� ܚ �� D� �� �� d� � џ �� @� �� �� i� #� ݤ �� R� � ɧ �� B� �� �� {� :� �� �� x� 9� �� �� ~� A� � ȳ �� P� � ۶ �� h� 0� �� �� �� R� � � �� }� I� � �� �� � N� � �� �� �� a� 4� � �� �� �� X� .� � �� �� �� d� =� � �� �� �� �� b� @� � �� �� �� �� �� b� E� (� � �� �� �� �� �� s� \� F� 0� � � �� �� �� �� �� �� �� }� o� a� U� I� >� 4� *� !� � � � �    �  � � � � � � � � �	 �
      # - 7 B N [ i w � � � � � � � ! "" :# R$ k% �& �' �( �) �* , 7- X. z/ �0 �1 �2 4 25 Z6 �7 �8 �9 ; 0< ^= �> �? �@  B SC �D �E �F *H cI �J �K M PN �O �P R OS �T �U W aX �Y �Z :\ �] �^ ` ma �b d `e �f h ^i �j l gm �n p }q �r <t �u w ex �y 2{ �| ~ o ܀ J� �� *� �� � �� �� s� � h� � b� � c� � i� � v� �� �� � �� 2� ä U� � � � �� J� � �� $� Ŵ i� � �� ]� � �� a� � �� v� +� �� �� V� � �� �� U� � �� �� s� ?� � �� �� �� ]� 5� � �� �� �� �� w� _� J� 6� %� � 	� �� � � � � �	 � � � 
  ' 9 N f � �  �" �$ ' )) S+ - �/ �1 4 M6 �8 �: = G? �A �C !F oH �J M mO �Q %T �V �X Q[ �] )` �b e �g �i }l �n �q 
t �v %y �{ M~ � �� $� Ȉ p� � ̐ � 6� � �� r� 9� � Ҧ �� {� U� 4� � �� � ڽ �� �� �� �� �� �� �� �� � -� N� u� �� �� � ?� ~� �� � Y� ��  c �	 / �  �  � " �% <) �, y0 !4 �7 �; <? �B �F �J bN ;R V Z �] �a �e �i �m �q v /z U~ �� �� � 5� �� ӗ .� �� �� m� � k� �� �� '� �� y� 0� �� �� �� d� I� 6� -� .� 9� N� l �	 �  M � �# d) �. V4 �9 t? E �J xP <V \ �a �g �m �s �y � � T� �� � K� �� 5� �� Z� � �� �� X� ?� 5� ;� R� z� �� � V � @ �# r+ '3 �: �B �J �R �Z �b :k �s �{ u� 	� �� u� M� <� C� b� �� �� Q� �� p� '� � � � # S- �7 ,B �L ~W Ub Lm cx �� � o� � ͱ �� �� �� ;� �� V�   *" o/ �< zJ AX 7f Zt �� 0� � ˮ � 2� �� o� `� �	 �	 �-	 f>	 ~O	 �`	 mr	 F�	 c�	 Ĩ	 k�	 [�	 ��	 �	 �
 
 x1
 :F
 Q[
 �p
 ��
 ��
 #�
  �
 ?�
 ��
 � ^) =B �[ Ju � ,� S� �� #� � 	7 �T &s � �� �� �� � 6 �X u| �� �� �� J �9 )b o� �� �� � +: nh ͗ R� � �, /a �� ��  �? I{ N� � v7 �y �  ZL ǖ x� �2 � D� */ �� �� �E �� � Hz �� <[ "� �M � �S �� �o � �� �I � �� �g �.  T�  ��! �" 
�# ��$ H�% $�& �( �a) W�* ^0, m�- [g/ n11 m3 �55 �y7 ��9 ߢ< 9�? >�B �xF �J �O �T ��Y �` �Lh �^q 7+| e=� �b� �֭ o�� �� �!��tX�	x:e`�/
Bad V_CopyRect Bad V_DrawPatch x=%i y=%i patch.width=%i patch.height=%i topoffset=%i leftoffset=%i Bad V_DrawPatchFlipped Bad V_DrawTLPatch Bad V_DrawAltTLPatch Bad V_DrawShadowedPatch TINTTAB XLATAB Bad V_DrawBlock pcx V_ScreenShot: Couldn't create a PCX   �?            ���            {�G�z�?CWILV%2.2d WIMINUS WILV%d%d WIURH0 WIURH1 WISPLAT WIA%d%.2d%.2d WINUM%d WIPCNT WIF WIENTER WIOSTK WIOSTS WISCRT2 WIOBJ WIOSTI WIFRGS WICOLON WITIME WISUCKS WIPAR WIKILRS WIVCTMS WIMSTT STPB%d WIBP%d WIMAP%d Could not place patch on level %d STFST01                                @�                                                           ��e     @�e     ��e             
   	                          �   �   �   �   E   z   �   f   t   Y   �   7   G   8   �      G      �      a   2   �   @   �   N   �   \   �   �   �   �   �   �   �   �   �   �   0   �   �   _   	  K   �   0        �   0   �        �                                                                           -mmap -file  couldn't open %s
 IWAD PWAD Wad file %s doesn't have IWAD or PWAD id
 Couldn't realloc lumpinfo W_GetNumForName: %s not found! W_LumpLength: %i >= numlumps W_ReadLump: %i >= numlumps W_ReadLump: only read %i of %i on lump %i W_CacheLumpNum: %i >= numlumps w_wad.c W_ReleaseLumpNum: %i >= numlumps doomgeneric 
You are trying to use a %s IWAD file with the %s%s binary.
This isn't going to work.
You probably want to use the %s%s binary. POSSA1 IMPXA1 ETTNA1 AGRDA1           B�C            I�C            P�C            W�C     Z_Free: freed a pointer without ZONEID Z_Malloc: failed on allocation of %i bytes Z_Malloc: an owner is required for purgable blocks zone size: %i  location: %p
 tag range: %i to %i
 block:%p    size:%7i    user:%p    tag:%3i
 ERROR: block size does not touch the next block ERROR: next block doesn't have proper back link ERROR: two consecutive free blocks ERROR: block size does not touch the next block
 ERROR: next block doesn't have proper back link
 ERROR: two consecutive free blocks
 Z_CheckHeap: block size does not touch the next block
 Z_CheckHeap: next block doesn't have proper back link
 Z_CheckHeap: two consecutive free blocks
 %s:%i: Z_ChangeTag: block without a ZONEID! %s:%i: Z_ChangeTag: an owner is required for purgable blocks Z_ChangeUser: Tried to change user for invalid block!                               	
 !"#$%&"()*+<_>?)!@#$%^&*(::<+>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[!]"_'ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~I_InitGraphics: framebuffer: x_res: %d, y_res: %d, x_virtual: %d, y_virtual: %d, bpp: %d
 I_InitGraphics: framebuffer: RGBA: %d%d%d%d, red_off: %d, green_off: %d, blue_off: %d, transp_off: %d
 I_InitGraphics: DOOM screen size: w x h: %d x %d
 -scaling I_InitGraphics: Scaling factor: %d
 I_InitGraphics: Auto-scaling factor: %d
 I_GetPaletteIndex LemonDOOM           zR x�  $      X0���   FJw� ?;*3$"       D   �2��-    Ak    \   54��           (   t   4��^    B�D�A �OAF     �   P4���    M�p     �   �4��1          �   �4���    A�   �   �5��J       (   �   �5��+   V�N�s ��AH     (  �6���          <  ^7��E   A?      X  �8��E    A�F |A    x  �8��6    A�F mA    �  �8��!          �  �8��u    As   �  ,9��&    Ad    �  :9��]    AW   �  9��#    A]      �9��#    A] (   $  �9��W   A�D�A NAA       P  �<��R    Ax
EI
EA (   t  �<���    e�A�A �AAA��    �  �=��N          �  �=��F    Jt
EA      �  �=��       8   �  �=���   B�B�A �A(�F0�(A ABB   0   $  �@��   h�N�P �G(�� ABB    X  {A��     A�X
EA ,   x  {A���    B�A�C �D0� AAB   �  B���    A��  8   �  �B��s    L�B�E �A(�D0�H(L BBB  D      "C���    B�E�E �E(�D0�C8�G`�8A0A(B BBBH   H  �C���    A�A�A n
(K0DH(K0H(B V(F0F(A RAA   4   �  XD��d    B�D�C �g(Z0I(E HAB   (   �  �D���    B�D�A ��AB     �  �D��%            E��t    Jd   $  kE��2          8  �E��2          L  �E��K    wJ    d  �E��#       H   x  �E���    B�B�D �D(�A0K
(A ABBEx(D ABB     �  BF��    A�P   H   �  8F���   B�B�J �B(�A0�A8�DP�8D0A(B BBB   4   ,  �G��k    B�J�A �C(�C0Q(A ABB   d  �G��%          x  �G��0          �  H��5              �  H��          �  H��?          �  6H��.    Al $   �  LH���    A�A�D0�CA(     �H��`    J�A�A PAAA��    8  &I���    D�c
E`   X  �I��    AS    p  �I��:          �  �I��     A�V   H   �  �I���   B�B�B �B(�A0�A8�A@�8A0A(B BBB      �  ?L��                /L��/            JL��K    \m    0  }L��0    K�d   (   L  �L��.   A�F�F0AA      x  �M��          �  �M��    AV @   �  �M��R   B�A�A �D0�
 AABEw AAB      �  �P���    A   �  XQ��          	  OQ���   A�      ,	  �R��       4   @	  �R���   A�A�A |
ICEAAA      x	  T���    A��     �	  �T��          �	  �T��)       ,   �	  �T��=	   B�I�A �A(�G�          �	  �]��'           
  �]��t          
  X^��-          (
  q^��3          <
  �^��          P
  �^��       8   d
  �^���    B�E�L �D(�D0��(A BBB     �
  _���    I`�   �
  �_��   D�  $   �
  �a��    A�K�A �AA8   �
  �b��   B�N�B �A(�A0��(A BBB     8  kc���          L  �c���   W�   $   h  Wg���    AZ
E^
EP      �  h���    vM   �  ph��       (   �  mh���    B�D�D ��AB     �  �h���    A�
EA     Ii��V       0     �i��_   B�K�A �D0H AAB      P  �j��x    `O       l  k��^          �  \k��       @   �  Kk��4   D�G�B �I(�G0�H8�0A(B BBB    �  ;l��          �  @l��)    Ag 4     Ql���    B�E�D �D(�A0f(A ABB(   <  �l���    D�D�L ��CB     h  Hm��%    Ac ,   �  Um��U    B�F�H �K0s CAB 8   �  zm���    B�E�D �C(�D0�(D ABB       �  �m��	       H      �m��Q   D�J�H �B(�A0�A8�D@(8A0A(B BBB      L  �s���   A�   (   h  Pu���   h�A�D {AA     �  x��V          �  Qx���          �  �x��       8   �  �x���   B�L�A �A(�A0�(A ABB   4     �z���    L�B�A �A(�C0s(A ABBd   D  �z���    V�B�B �A(�R0�U
�(A� B�B�B�EQ
(I BBBAJ�(D� B�B�B�   �  F{��          �  ={��          �  >{��A    J`    �  g{��}   Au
A     �}��`             ~��4    Ar    8  ,~��    A]    P  3~��"    A` (   h  =~��7   B�A�A �AB    �  H��       8   �  Q���   B�B�D �C(�C0�(A ABB   $   �  ����    A�D
Ee
EA      �����    A�$   $  ����    A�J�A �AA   L  ����?    kR    d  ����U   AS      �  ����       (   �  ����   B�M�A ��AR    �  ����;    A�U      �  ܅��X   AV      �  ����       L     ����D   I�B�J �D(�A0��
(A BBBEd(D BBB   �   \  ����;   B�B�A �A(�D0�
(A ABBEP
(A ABBEA
(A ABBEA
(A ABBEA(A ABB          �  5���          �  "���             ���             +���*          4  A���#       H   H  P����    B�B�E �D(�A0��
(A BBBEA(A BBB4   �  �����    B�B�A �A(�D0�(A ABB   �  '���l          �  ���Z          �  Ō��V       $     ���D    N�D�C lAA $   0  #���U    A�C�D JAA   X  P���4          l  p���          �  j���          �  l���          �  q���#          �  ����?    A�}      �  ����          �  ����3    A�q            ����F    A�F }A    ,  ܍��       4   @  Ӎ���   A�A�A [(M0�(A �AA      x  J���-    Ae
EA      �  W���     AZ 8   �  _����   H�B�B �A(�A0��(A BBB    �  ݐ��6             ����%       ,     ����   A�A�A zAA          D  `���              \  I���          p  6���          �  #���       (   �  ����    A�P�F@�AA    (   �  ����y    B�F�A �lAB     �  ���8    MT
BA        ���          $  ����B    MY
BA      D  !���5          X  B���>          l  l���          �  h���          �  f���          �  j���          �  W���          �  D���          �  @���          �  <���            8���             6���          4  2���          H  .���          \  *���          p  (���       $   �  ���.    A�I�C ^AA    �  ���       (   �  ���E    B�J�F �kAB      �  !���    A�Y        $���-    D g       9���          4  (���    A�U   (   P  #���8   B�B�A �D(�G�   (   |  /���u    B�F�I �`AB  H   �  x����   B�B�E �B(�A0�D8�FPp8A0A(B BBB      �  ����            ����+    Ai       ×��    A]    8  ʗ��          L  ����          `  ����       8   t  ����K    B�E�I �A(�G0�h(D BBB      �  ����          �  ����    AF    �  ����          �  y���&    H�]        ����             ����"          4  �����          H  ���       8   \  ���F    B�E�B �D(�C0�n(A BBB   $   �  ���F    A�L�A uAA    �  8���9    D t    �  Y���          �  T���             A���            .����    A�
E_     4  ˘��    A�T   $   P  Ř���    A�D�A �AA   x  2���#    Aa    �  =���%    Ac    �  J���$    Ab    �  V���J    AD   �  ����D    W�l      �  �����   A�        +����    A�   (  �����    A�   @  +���.   A(      \  =����    A�   t  �����    A�   �  ����y   As   $   �  ����Q    A�M�F@zAA    �  ���          �  
���          �  ���:            .���K             e���'    A^    8  t���#    AZ    P  ���D    A{    h  ����#    AZ    �  ����6    G�n$   �  Ԡ��i    A�A�A cAA$   �  ����    A�A�A �AA   �  ����7          �  ء��7            ����U    AS   (  8���R          <  v���+          P  ����S    Ry    h  Ȣ��"    IS    �  Ң��.    Ic    �  ���*       0   �  �����    B�A�F �I�� AAB   (   �  v���p    B�A�H �ZDB        ����4    D�o      (   ң��"    IS D   @   ܣ���    B�B�E �E(�I0�C8�I@�8A0A(B BBB   �   L���f    A]   �   �����    A�$   �   U���4    A�I�H QHD $   �   a���4    A�I�H QHD    !  m���5          !  ����a    oh    4!  ץ��=          H!   ���Y    FI   `!  A���9    Z^    x!  b���       (   �!  e���Q    B�G�C �AAB     �!  ����:       8   �!  ����n    B�E�E �D(�C0�S(A BBB  $   "  ���h    A�P�C QAA0   0"  "����    A�K�C �
EAEAAA   d"  ����,       @   x"  �����   B�B�B �A(�A0�D��0A(A BBB     �"  g���          �"  ^���          �"  \���(    XK    �"  l���2    aK    #  �����    _j
Al   (   4#  ���	   I�A�D �	AB    `#  Բ��
          t#  ʲ��A          �#  ����Q    AK   �#  0���
          �#  &���
          �#  ���
          �#  ���!          �#  ���'          $  2����              $  ֳ��
          0$  ̳��>    A| (   H$  ���>    B�A�A �vAB   (   t$  ���H    B�I�C �vAB   D   �$   ����    B�B�J �B(�D0�A8�A@p8A0A(B BBB$   �$  i���m    A�I�I WAA4   %  ����u    B�J�D �V
CBEAAB     H%  ���    A�Y   D   d%  ���t    B�H�B �E(�D0�A8�A@O8D0A(B BBB$   �%  ���9    A�A�D pAA    �%  '���>    I�kG� D   �%  I���   B�G�E �F(�D0�G8�DP�8D0A(B BBB   8&  ���$          L&  ���A    lI    d&  ;���B    iM 0   |&  e���$   B�F�A �Dp DAB      �&  U���       (   �&  W���/    H�D�E ZAAA��     �&  Z����    G��      '  ȷ��           '  ͷ��          4'  ҷ��              L'  Ϸ��"          `'  ݷ��:    A�x   4   |'  ����H   A�A�D w
DAE�AA      �'  ���6       H   �'  -���&   E�B�E �B(�D0�A8�A@8C0A(B BBB      (  ���B           4   ,(  1����   J�i�c��
�EY
�EAA�   H   d(  ����u   B�L�E �E(�E0�A8�C@G8C0A(B BBB      �(  Ӽ���    h�
AA  ,   �(  m���"   ��D�A �pABA���$    )  _���R    A�K�F }AA (   ()  ����n    A�K�F YAA       T)  ˿���    jf<   l)  K����    Y�E�A �C(�D0�(A ABBA����      �)  ����       $   �)  ����V    A�A�A PAA$   �)  ����   A�D�A �AA(   *  ����   B�A�A �AB    <*  ����"    A�`   H   X*  ����D   B�B�B �B(�A0�A8�GP(8A0A(B BBB   D   �*  ����   B�B�H �E(�A0�A8�GP�8A0A(B BBB   �*  ����b    FpZ   +  �����    A��
HA,   $+  v����   A��
E}
E�
HA   (   T+  =���V    M�A�D @AAA�� 8   �+  g���    L�B�A �A(�D0F(H� H�B�B�L   �+  �����    P�M�B �B(�G0�A8�D@_8A0A(B BBBA������ 8   ,  ����    L�G�A �A(�D0A(H� H�B�B�   H,  5���I    A�i
HV    h,  ^���I    A�i
HV    �,  ����)    K�S�      �,  ����g    K�A
�EP�      �,  ����I    K�v
�EAA�      �,  ����Z    K�t
�EP�      -  2���)    K�S�      ,-  ?���_    K�y
�EP�      P-  z���R    K�EA�,   l-  ����`   O�A�A �JABA���    �-  ����"    K�Q�  (   �-  ����h    K�G ~
L�EDAA� `   �-  "���e   B�B�B �B(�A0�D8�A@)
8A0A(B BBBAQ8D0A(B BBB      H.  #���
       H   \.  ����    B�B�A �A(�A0�
(A ABBEA(A ABB     �.  g���    A�Q      �.  b���    A�Q      �.  ]���R    K�A� P   �.  �����    P�B�A �A(�D0�
(A� A�B�B�EA(A ABBA����    P/  ,���    A�Q   $   l/  '����    A�A�D �AA$   �/  �����    A�A�D �AA4   �/  �����    B�B�D �A(�A0�(A ABB(   �/  �����    B�A�A ��AB  T    0  "����    w�M�B �D(�C0��
�(A� B�B�B�ES�(A� B�B�B�     x0  ����     K�O�     �0  ����<    A�p      �0  ����`    A�X
EA   �0  +���
          �0  !���          �0  !���          1  ���           1  ����   (p{     <1  ����    A�Q      X1  ����    A�Q      t1  ����    A�Q      �1  ����          �1  ����       $   �1  ~���$    A�I�D IGA    �1  z���e          �1  ����       4   2  �����    B�E�A �F(�A0�(F CBB(   @2  1����    B�A�D �uAB     l2  ����       (   �2  v����    _�A�D [A�A�  (   �2  ����   M�D�A �D�A�     �2  ����    A�Q      �2  ����#           (   3  ����	   B�A�C ��AB  0   83  �����    A�D�D |
AAIAAAH   l3  ����W   B�G�B �H(�D0�A8�DP.8C0A(B BBB   H   �3  �����   B�E�E �E(�D0�D8�D`r8D0A(B BBB   ,   4  L���1   K�D�C �ABA��� 4   44  M���   B�B�A �C(�G0�(D ABB   l4  ���)          �4  .���          �4  0���          �4  :���x       <   �4  ����R   i�D�A �
�E�B�EAABA���     �4  �����   A�� �   5  I���   P�B�B �B(�A0�A8�GP
8G�0A�(B� B�B�B�E�
8D�0A�(B� B�B�B�ER8A0A(B BBBA������          �5  ����+          �5  ����M          �5  ���:    F�rA�    �5  &���=    M�nA� $   6  G���T    A�K�A DAA$   46  s���d    A�K�A TAA4   \6  �����    B�J�F �I(�A0g(A ABB$   �6  ���@    A�D�D tAA 8   �6  ���n    B�E�E �A(�A0�X(A BBB  8   �6  K���p    B�E�E �A(�C0�X(A BBB  $   47  ���U    A�K�F @AA    \7  �����   A�I �C   $   �7  L����    A�D�A �AA8   �7  ����e   B�B�D �A(�A0R(C ABB   H   �7  �����   B�B�B �B(�A0�D8�A@�8D0A(B BBB      08  l���|    aS   H8  �����   }�sA�      h8  g���e    A�c  (   �8  �����    \�A�A gFAA�� H   �8  ���p   B�G�E �B(�A0�A8�DPO8A0A(B BBB   8   �8  ;����   B�D�B �A(�A0��(A BBB H   89  ����e   B�B�E �B(�A0�C8�D@G8A0A(B BBB   (   �9  ����X    B�A�A �JDB  $   �9  �����    A�A�D �FA(   �9  �����    j�A�A ��AH  `   :  ;����   B�B�H �H(�A0�A8�GPu
8A0A(B BBBE�8A0A(B BBB   $   h:  �����    A�C�C �AA   �:  C���z          �:  ����G       8   �:  �����    B�J�L �A(�A0�g(A BBB  ,   �:  )���L    R�A�D �kGB          $;  E���t          8;  ����1          L;  ����#       ,   `;  ����m    w�G�C �^AEG���   (   �;  ����    B�A�A ��AB  ,   �;  �����    C�C�C �|ABA���     �;  
���       H    <  ���s    B�E�A �A(�E0J
(C EBBEA(C ABB  $   L<  7���
   A�A�G0�CAD   t<  ����    B�B�B �E(�A0�A8�D`�8F0A(B BBB   �<  ����Y          �<  �����          �<  �����    A��  (    =   ���}    ^�D�A QAAA�� (   ,=  q���W    ^�D�A kAAA��  4   X=  ����s    B�E�D �C(�A0](A ABB`   �=  ����b   B�E�E �B(�A0�A8�Dp)
8F0A(B BBBED8C0A(B BBB   8   �=  � ��+   B�J�J �D(�E0�(A BBB    0>  ����    A��  $   L>  6��z    A�A�D qAA   t>  ���m    A�e
EA4   �>  ����   A�A�D 
DAE^AA  T   �>  #��5   z�B�B �A(�A0��
�(A� B�B�B�E�(A BBBA�����4   $?   ��   B�A�A � 
ABEAAB $   \?  ����    A�j
H~
EA  <   �?  i��2   O�B�A �A(�A0(A ABBA����  <   �?  [��L   Q�A�A �+
�A�B�EAABA���  ,   @  g	���   ��C�D !AAA��   0   4@  ���    A�C�D0j
IAEDAA<   h@  h���    B�D�C �D0y
 AABED AAB    �@  ���[    A�S
EA   �@  ���-       8   �@  ��   B�D�E �A(�D0��(A BBB  8   A  ���   B�J�B �D(�A0��(A BBB     TA  ���2          hA  ���<          |A  ���-       H   �A  ���   B�E�E �B(�A0�D8�DP�8C0A(B BBB      �A  ���E    A�m
AQ D   �A  ���.   A�A�D �
DAEZ
AAEAAA          DB  ���       4   XB  ����    B�E�A �D(�E0�(A ABB   �B  +��M    AK   �B  `��[    A�U     �B  ���_   }       �B  ���?    A�t
HA     C  ��       @   C  ��    B�D�A �\
ABOh
ABEMAL    XC  ���/          lC  ���          �C  ���>          �C  ���.          �C  ��,    A�\   ,   �C  ���    B�A�D �D0� AABH   �C  ����    B�B�A �D(�A0j
(A ABBEu(A ABB    @D  K��&    A`    XD  Y��&    A` $   pD  g��R    A�F�D @AA$   �D  ���e    A�D�A \AA,   �D  ���e    B�D�A �F0E FFB   �D  ��m    A�g  $   E  T��p    A�K�D ]AAD   4E  ����    B�G�H �H(�A0�A8�D@�8A0A(B BBB0   |E  0���    A�I�D �
AAEAAA   �E  ���          �E  ���          �E  ���       4   �E  ����    B�B�A �D(�C0�(A ABB   $F  ���          8F  ���$       $   LF  ��[    A�C�D PAA   tF  4��R    D M   �F  n��    A�O      �F  d��-    A�g      �F  u��    A�W      �F  s��^    A�X  $   �F  ���+    A�C�A cAA    $G  ���Q    D L   <G  ���    A�V   (   XG  ���7    B�A�A �jFB   $   �G  ���)    A�C�A aAA    �G  ���&    A�d      �G  ��8    Kd    �G  #���    A�F0{A,    H  ����    B�D�A �F0� AAB,   0H  0���    B�A�A �I@� CAB   `H  ���    AF    xH  ���
       8   �H  ����   B�L�B �G(�A0��(A BBB 8   �H  =���   B�B�G �A(�C0�(A ABB   4   I  ����    B�B�A �C(�A0�(A ABB4   <I  w ��	   B�B�A �C(�A0�(A ABB(   tI  H!���   A�K�A �CA      �I  #���   A��    �I  �%��d   A�H
E     �I  �'���   A��        �I  f+��p    A�j     J  �+��W    T| 8   0J  �+��C   B�E�A �C(�A0*(C ABB      lJ   -���    A��  4   �J  p-���    B�E�D �A(�A0�(D ABB   �J  .���    A��  4   �J  �.���    B�G�D �C(�D@�(A ABBH   K  3/���   B�B�B �E(�D0�A8�A@p8D0A(B BBB   4   `K  z0���    B�E�A �C(�A0�(C ABB   �K  $1���    A��  8   �K  �1��?   B�D�A �A(�D@,(A ABB   8   �K  �3���   B�I�E �A(�F`�(A ABB      ,L  +6��    AP    DL  )6��h       H   XL  }6��s    B�E�A �A(�E0J
(C EBBEA(C ABB  H   �L  �6���   B�B�B �B(�A0�A8�G`�8A0A(B BBB   4   �L  08���    [�A�A u
A�A�EFAA     (M  �8���       4   <M  T9���    B�B�A �A(�F0�(A ABB   tM  :��.          �M  :��2          �M  ::��!          �M  G:��          �M  I:��4          �M  i:��7       H   �M  �:���    B�E�B �E(�D0�C8�F�q8C0A(B BBB      8N  �:��8          LN  �:��5          `N  ;��4          tN  >;��6       X   �N  `;��F   A�b
E�
EJ
ED
EP
ET
E|
E`
EI
EP
EA     �N  J>��k    A�c
EA,   O  �>���    A�d
E\
EH
EA   (   4O  ??��_   I�A�A �PAB H   `O  r@��$   B�E�B �B(�E0�A8�DP8D0A(B BBB   ,   �O  JB���   A�A�A �AA       8   �O  �C���    B�B�G �A(�A0G
(A ABBA    P  D��~       4   ,P  �D��Z   B�D�D �@
DBEAAB    dP  �E���   ]�KA�  <   �P  5H���   D�B�B �A(�A0�@(A BBB       �P  �I��          �P  �I��          �P  �I��	           Q  �I��          Q  vI��E    A�C     0Q  �I��x    Q�eA�(   LQ  �I��B    L�D�F �hAB   $   xQ  J���    A�A�D �AA   �Q  �J���    A�~
EA   �Q  NK���    A��     �Q  �K���   @��       �Q  �M��       (   R  �M���    B�G�C ��AB  0   <R  |N��Y    A�F�F 
CAEAAA    pR  �N��-       <   �R  �N��   A�D�A �
CAEA
CAEAAA,   �R  �O��"   }�E�O ��CBA���  $   �R  ~P���    A�A�D �AA4   S  .Q���    [�A�A e
A�A�BAAA     TS  �Q��N       D   hS  �Q��   B�G�B �B(�A0�A8�GP�8N0F(B BBBH   �S  �R���   B�M�E �B(�A0�I8�DPY8A0A(B BBB   $   �S  �S��n    A�D�A eAAH   $T  T��   B�L�B �B(�A0�C8�D��8A0A(B BBB     pT  �X��b    A`$   �T  #Y���    A�F�C �AA   �T  �Y��     A^    �T  �Y��1    An $   �T  Z��B    A�D�D0vAA (   U  *Z��T    H�D�A CAAA�� $   4U  RZ��&    A�D�A ]AA L   \U  PZ��}   O�G�B �B(�A0�A8�A@M8D�0A�(B� B�B�B�    �U  }\���    M��     �U  ]���    M��     �U  �]���    H��  (    V  �^��   A�A�A AA      ,V  p_���    M��  $   HV  `���    A�A�A �AA   pV  �`���    A�   �V  Va���    A�   �V  b��   A      �V  c��f       4   �V  Sc��q   A�A�A c
AAEAAA      W  �e��%          W  �e���    X�   4W  2f��       ,   HW  =f���    C�C�C �tABA���  ,   xW  �f���    l�A�A �QABA���     �W  �f��   g�   �W  �g��          �W  �g��e    O�y      �W   h��       $   X  h���    F�A�C {AA   ,X  mh��       (   @X  Zh��   N�D�D ��AB  4   lX  =i���    B�H�D �A(�F0k(A ABB   �X  �i��       (   �X  �i���   A�A�A |AA      �X  �k���    A�(   �X  Ql��]    T�G�C �nAD      (Y  �l���          <Y  -m��G    AA   TY  \m��       H   hY  Im���   B�B�B �E(�D0�C8�DPi8A0A(B BBB      �Y  �n���    M��  4   �Y  o���    B�G�D �C(�F0z(D ABB   Z  io��       D   Z  �o���    B�E�E �E(�D0�D8�GP�8A0A(B BBB<   dZ  ?p��   I�B�I �A(�A0��(A BBB     8   �Z  r��   B�B�A �C(�A0(A ABB   8   �Z  �s��   B�B�B �A(�D0��(A BBB L   [  �v��{   S�B�B �B(�D0�A8�FPK8A0A(B BBBA������   l[  �~��           H   �[  �~��B   B�B�E �E(�D0�C8�B@ 8A0A(B BBB   L   �[  ���Z   f�I�B �B(�A0�F8�I`8A0A(B BBBA������    \  ���          4\  ���          H\  ���!       $   \\  ����    A�A�D �AA8   �\  ����!   B�G�A �A(�D0(A ABB   H   �\  w����   B�E�B �B(�A0�A8�DP�8A0A(B BBB      ]  ͅ��j    L�\A�H   (]  ����   B�B�B �E(�A0�A8�D��8A0A(B BBB     t]  �����    A��
EA   �]  +����       8   �]  ���   B�B�D �A(�A0�(A ABB      �]  Њ��q    A�i
EAH   ^  !���+   B�F�B �B(�A0�A8�DP8A0A(B BBB      P^   ���,       8   d^  ����    B�B�B �D(�D0��(A BBB  4   �^  �����    B�B�D �A(�F0�(A ABB   �^  ���    D Y    �^  ����          _  ����D    A�B      _  ����          4_  ����    AW    L_  ����        l   `_  ����A   B�B�B �B(�A0�D8�DP�XN`LXAPo
8E0A(B BBBED8A0A(B BBB      �_  ����          �_  {���#       $   �_  ����-    A�C�D \FA     `  ����       H   4`  �����    m�B�A �A(�G@HHNPOHA@f(A ABBA����      �`  ���       \   �`  ����    b�B�B �B(�A0�A8�E@OHLPVHA@J8A0A(B BBBA������        �`  p���    A�Q   @   a  g���`   B�B�B �A(�C0�G@F0A(A BBB      Ta  ����    A�P      pa  y���q    JIS I  ,   �a  ʡ���   B�A�G0[CAA��      �a  G���A          �a  t����   A�      �a  <����    A�   b  
���)    Ag     b  ����    H��
EA$   @b  �����    A�C�C �HA   hb  ����    AU    �b  ����          �b  {���A    Fv
BA      �b  ����
          �b  ����    AQ    �b  ����
          �b  ����          c  r����       L   c  ����   I�L�Q �F(K0a(^0}(B O(Q0|(P00(A AAB   lc  6���/    Jc    �c  M���%    Ac    �c  Z���     A^    �c  b���    AF    �c  V���8    A�v   8   �c  r���   B�E�A �A(�B0(A ABB      $d  J���/       8   8d  e����   B�B�D �A(�G@�(A ABB      td  ����&    TP    �d  ���&    TP <   �d  ����    B�B�B �D(�A0�F@�0A(A BBB   �d  ����    A�X       e  ����    A�\   $   e  �����    A�H�H wFF   De  ���          Xe   ���Z    KM$   pe  B����    A�C�D0�AA   �e  ݳ���    A�F@rF   �e  A���          �e  4���)           8   �e  E���K    R�E�F �E(�H0F(P� A�B�B� D    f  T����    B�E�E �E(�D0�C8�DP�8A0A(B BBB   hf  ���       4   |f  ش��   B�A�D �[(T0H(A AB (   �f  �����    B�A�D ��AB     �f  l���       (   �f  ]����    B�A�D ��AB  (    g  ����    B�A�D ��AB  (   Lg  �����    B�A�D ��AB  D   xg  <����    B�B�B �B(�D0�A8�A@�8A0A(B BBB   �g  ���    AW    �g  ���    AW 8   �g  ����    B�E�E �D(�D0�o(A BBB     ,h  B���:          @h  h���%          Th  y���,          hh  ����:    A�w      �h  ����          �h  ����          �h  ����          �h  ����       D   �h  ����   B�E�E �N(�F0�D8�LP�8D0A(B BBB$   i  N���v    A�D�F0hAAd   Di  �����   B�L�B �B(�A0�A8�KPm
8I0F(G BBBED8A0A(B BBB          �i  ���    A�Q   H   �i  ���@   B�B�B �B(�A0�C8�G`"8A0A(B BBB      j  ۾��    A�P      0j  Ѿ��          Dj  ;��       $   Xj  �����    A�A�DP�AA$   �j  Q���n    A�F�F XAA   �j  �����       ,   �j  F����    _�A�C �{ABA���  ,   �j  �����    _�D�A ��ABA���     k  h���W    V�A� D   8k  �����    B�E�E �B(�D0�C8�DP�8C0A(B BBB(   �k  /���/    F�K�C �R�A�B�T   �k  2����    J�B�E �D(�C0�m
�(A� B�E�B�GA(A BBBA�����    l  z���          l  ����    AN
EA      8l  {���#          Ll  ����6    A_
BS   0   ll  �����    A�A�A o
AAEkAA   �l  ���          �l  ���2          �l  ,���t       $   �l  �����   A��
EA
E_ H   m  N����   B�B�B �B(�A0�F8�C@�8A0A(B BBB      Pm  �����    A�$   hm  c���    A�
EA
E_   H   �m  [���9   B�B�B �B(�A0�A8�F@8A0A(B BBB      �m  H���_       $   �m  �����   A`
EA
E_   0   n  ����   A�F�A �
FAEAAA   Ln  �����       4   `n  R���|    BH
EK
EJ
EA
EA
EA     �n  ����r    Ap   �n  ����
          �n  ����          �n  ����?          �n  ����v            o  a���/    AT
EJ
EA L   $o  l���   B�B�B �B(�A0�C8�G��8A0A(B BBB          to  ���    A�X      �o  ���          �o  ���           ,   �o  ����k    B�K�A �YAB      (   �o  8���6    B�D�C �iAB   H   p  B���\   B�B�B �B(�A0�A8�G`=8D0A(B BBB      dp  R���       (   xp  E����    B�D�H ��AB  $   �p  ����&    A�D�A ]AA    �p  ����)    A�g   (   �p  ����f    H�D�C �MCB  4   q  �����    B�E�D �A(�A0�(D ABB   Lq  W���    D Q    dq  [���K    A�~
JA    �q  ����    AF 4   �q  y����    B�B�A �A(�A0(A ABB4   �q  �����    B�B�D �A(�F@l(A ABB   r  ���7           r  ;���T    D O$   8r  w����    A�E�D �AAD   `r  ����   B�H�E �E(�E0�A8�A@�8A0A(B BBB(   �r  ����P    I�A�C �AB   (   �r  �����    I�D�H ��AB  $    s  z����    A�I�A �AA   (s  ���q    H�h  4   Ds  Y���V    B�E�D �C(�E0|(A ABB $   |s  w���*    A�D�D ^AA    �s  y���,          �s  ����
       (   �s  ����2    B�F�F �TIB      �s  ����    A�P   $   t  ����P    A�F�A EAA   <t  �����    D0�   Tt  F���              lt  /���a          �t  |����    P��  $   �t  +����   Z�M G(G0K�   �t  ����    AT    �t  ����          �t  ����          u  ����       D   u  u����    B�B�B �B(�A0�A8�A@�8A0A(B BBB   `u  ���          tu  ����]       (   �u  G���I    B�D�G �xAB      �u  d���          �u  Q���          �u  >���          �u  /���          v  ���          v  	���          ,v  ����          @v  ����          Tv  ����              lv  ����    AT    �v  �����    A��     �v  L���E    AC   �v  y����    D@   �v  ����    C�T      �v  ����&    A�d      w  ����2          w  	���$    A�\
EA    <w  ���              Tw  ����1    A�CA�k   tw  ���D    A�CA�~   �w  *���8    A�Cs      �w  B����    A�C�     �w  �����    A�C�     �w  ����u    A�Cp      x  ����[    A�CA�U      8x  ���.    A�Ci      Xx  )���I    A�CD     xx  R���   A�C    �x  J���Q    A�CL     �x  {���J   A�CE    �x  ����j   A�Ce    �x  ����W    A�CR     y  &����   A�C�    8y  �����    A�C�     Xy  L���?   A�C:     xy  k���    A�C        �y  g���>    A�CA�x   �y  ����D    A�CA�~   �y  ����/    A�CA�i   �y  ����0    A�CA�j   z  ����2    A�Cm      <z  �����    A�C{      \z  ����   A�CE��      �z  *���    A�CV      �z  F���C    A�CE�y   �z  i���6    A�CA�p   �z  ����    A�C}      {  �����    A�C�      {  �����    A�C�     @{  #���    A�Cz     `{  �����    A�C�     �{  R���&    A�Ca      �{  &���-    A�Ch      �{  4���-    A�Ch      �{  B���    A�CL       |  4����    A�C�      |  ����"    A�C]      @|  ����"    A�C]       `|  �����    A�CE��      �|  J���-   A�C(    �|  $���)    A�Cd      �|  -���)    A�Cd      �|  6���    A�CV      }  1���    A�CZ      $}  0���    A�CV      D}  +���    A�CZ           @     ��������        ��������                             0@            �JB            0Yd                          h@            �@            �@     
       6                                          �Zd            �                           X@            (@            0       	                                                                                                                      XYd                     V@     f@     v@     �@     �@     �@     �@     �@     �@     �@     �@     @     @     &@     6@     F@     V@     f@     v@     �@     �@     �@     �@     �@     �@     �@     �@     @     @     &@     6@     F@     V@     f@     v@     �@     �@     �@     �@     �@     �@     ��������                xma                        ema                                       iddt                                                                      33                   ����L��               ���3�   ���3�   ����L��                "�� �����   �����   ���              "�� ���                  ��    $I     $I     �$	 0 $I     �$	 ����  ��    �m��0   ��    �m������I���      ��0 I���      ������n���    n�������n���������������������������I� ����    ����������������    ����    ����    I� 0 I� 0 Dc��0 Dc��y� ����y� ����M� Dc��  ��    $I     $I     �$	 I� $I     �$	 �m��  ��    �m��I�   ��    �m���m��I���      ��I� I���      ���m��              �KB     �KB     �KB     *LB     ^LB     �LB     �LB     
MB     �KB     EMB     wMB     �MB     �MB     NB     MNB     �NB                                  
                               3   2   1   4   7      ;   :   9   <   ?      L   K   J   M   O      S   R   Q   T   X      F   E   C   G          "   !       #   /      ����                              y0@     �W@     �D@     ۲@     aB            aB            +aB     
       =aB            OaB            AaB            KaB            UaB            aaB            oaB            {aB            �aB            �aB            �aB            �aB            �aB            �aB                                           �aB     �aB                   �cB     �cB                   qeB     yeB                   fgB     ngB                  fiB     niB                  kB     kB                  vmB     ~mB                  �nB     �nB                  �pB     �pB                  [qB     cqB                  fiB     �qB                  kB     FsB                  vmB     }tB                  �nB     �uB                  �pB     5wB                  [qB     �wB                  fiB     EyB                  kB     �zB                  vmB     �{B                  �nB     }B                  �pB     �~B                  [qB     oB        Z   x   x   Z   �   x   x     Z   �   �   �   �   �   �   �  �   �   �   �   �   �   �   �   ,  J  �  ,  �   x                                                     K   x   Z   �   �   �      �       Z   Z   Z   x   Z   h  �      �       Z   -   Z   �   Z   Z   �      �         �     @         (      2                          H�B     Z�B     n�B     ��B     ��B     ��B     ƅB     ۅB     ��B     �B     �B     =�B     S�B     f�B     ��B     ��B     ��B     ��B     ؆B     �B      �B     �B     *�B     C�B     W�B     l�B     ��B     ��B     ��B     ևB     �B     �B     �B     "�B     9�B     H�B     W�B     k�B     ��B     ��B     ��B     ��B     ˈB     ܈B     �B      �B     �B     )�B     <�B     O�B     e�B     s�B     ��B     ��B     ��B     ЉB     �B     �B     �B     5�B     J�B     f�B     ��B     ��B     ��B     ��B     ԊB     �B     ��B     �B     "�B     2�B     A�B     U�B     j�B     ��B     ��B     ��B     ȋB     ܋B     ��B     �B     �B     =�B     Z�B     z�B     ��B     ��B     ��B     ҌB     �B     ��B     
�B     �B     3�B     E�B     Y�B     f�B     z�B     ��B     ��B     ��B     ύB     �B     ��B     �B     $�B     ;�B     J�B     [�B     p�B     ��B     ��B     ��B     ͎B     ݎB     ��B     �B     �B     2�B     C�B     O�B     Y�B     g�B     z�B     ��B     ��B     ��B     ϏB     �B     �B     �B     #�B     #�B     #�B     #�B     #�B     #�B     #�B     #�B     #�B                             ,�B     4�B     =�B     E�B     K�B     N�B     f�B     n�B     ��B     ��B     ��B     ��B     ��B     ϐB                     �����   d   �               �   �          �   �   �   9            8 d                �  �      �   $         �   �          �   �   �   ;           8 d       K    @ �   	   �      �   %          �   �          �   �   �   <           8 d       K    @ �   @   �   �  �   0            
          �         G           8 �      P    @     ����  �                                                           d                 B   A  ,  C  j          W  d      O  S  Y      J   
        8 �      i    @ _  ����<  �      k                              >      R     
       d   
            ����7  �                                                           d                 C   j  X  l  1          �  P          x  �      d        0   @ �      K    @ �  ����e  �                                    g                  d               A   �  F   �  %          �  �          �  �  �  <           8 d       K    @ �  �  �  <   �  '          �  �      �  �  �  �  >           8 d       L    @ �  �  �  �   �  )      4   �  �      �      �      @   
        8 �      M    @ �  :   �  �   �  )      4   �  �      �      �      @   
        8 �      M    D �  �  �  �  �  *          �  �          �  �      A           8 �      M   B@   �    �    +            2                C           @ �      M    @ %  ����
  �                                                      d               E   ,  �  .  /          9  2      6  6  ;      H           @ �      M    @ B  �  I  d   K         3   Q            M  S                 8 2      M   B         Y  �  [  -         k  (          g  m      E        �   d �      M    @     D   x  �  z  .          �  �          �  �      F        @   @ X      N    @ �     �  �  �  ,          �            �  �      D        (   n �      M    @     G   �  �  �  2          �  �          �  �      I           8 �      M   B@ �  T   �  2   �  e          �  �          �  �  �  f           8 d       K    @ �  H   �  d                       g           �      h            H ���         @     X   
  �                    �   a                 b             ���                Y     �                                                          d                  W       �                                                            d                  ����  �      ^                                           
        d               ����  �                                                           d                 �  &                                        (      R         
   * d                 ����a   �                                    c            
       d               ����f   �                                    h            
       d               ����r   �                                           R            d               ����k   �                                    m                   d               ����s   �                                     u                   d   d            �����  �                                    �                  d               ����]   �                                                           d                 ����Z   �                                                           d                  �����   �                                                           d                 �����   �                                                           d                        �                                                           d                  ����{   �                                                           d                 �  "  �                                                           d                  �  $  �                                                           d                  �  0  �                                                           d            �     �  6  �                                                           d            �        <  �                                                           d                    >  �                                                           d                    @  �                                                           d                 '   F  �                                                           d                 &   D  �                                                           d                 (   B  �                                                           d                 �  H  �                                                           d                  �  I  �                                                           d                  �  J  �                                                           d            �     �  P  �                                                           d            �     �  T  �                                                           d            �     �  U  �                                                           d            �     �  ]  �                                                           d                  �  ^  �                                                           d            �     �  d  �                                                           d            �     S   Y  �                                                           d            �     �  f  �                                                           d                     g  �                                                           d                  �  h  �                                                           d                  �  i  �                                                           d                  �  j  �                                                           d                     k  �                                                           d                  �  l  �                                                           d                    m  �                                                           d                     n  �                                                           d                  �  o  �                                                           d                  �  p  �                                                           d                  �  q  �                                                           d                  �  r  �                                                           d                  �  s  �                                                           d                  �  t  �                                                           d                  R   u  �                                                           d                  U   �  �                                                           d                  V   �  �                                                           d                  �  v  �                                                           d                     �  �                                                           d                     �  �                                                           d                      �  �                                                           d                  !   �  �                                                           d                  %   �  �                                                           d                  $   �  �                                                           d                  )   �  �                                                           d                  *   �  �                                                           d                  +   �  �                                                           d                  ,   �  �                                                           d                  -   �  �                                                           d                  .   �  �                                                           d                  7   �  �                                                           d                  8   �  �                                                           d                  9   �  �                                                           d                  /   �  �                                                           d                  0   �  �                                                           d                  "   �  �                                                           d                   #   �  �                                                           d                  1   x  �                                                          D d                 2   �  �                                                          T d                 3   �  �                                                          T d                 4   �  �                                                          D d                 5   �  �                                                          4 d                 ;   �  �                                                          T d                  <   �  �                                                          D d                  =   �  �                                                          4 d                  >   �  �                                                          4 d                  ?   x  �                                                          D d                       �                                                           d                      �   �                                                           d                      �   �                                                           d                      �  �                                                           d                      X  �                                                           d                      �  �                                                           d                      �   �                                                           d                   
   �   �                                                           d                      �   �                                                           d                      ~  �                                                           d                       �                                                           d                      �  �                                                           d                     �  �                                                           d                     �  �                                                           d                     �  �                                                           d                  6   �  �                                                            d                  F   -  �                                                           d                  I   �  �                                                          X d                 J   �  �                                                          X d                 K   �  �                                                          @ d                 L   �  �                                                          @ d                 M   �  �                                                          @ d                 N   �  �                                                          @ d                 O   �  �                                                           d                  P   �  �                                                           d                  Q   �  �                                                           d                              ����                                          -9A                                   �1A                                  3A                                  S3A                                                                     �3A                                                                             	                            �2A                                  �1A     
                             3A                                  S3A                                                                      �6A                                                                     �2A     
                   �         89A                                  �1A                                  3A                                  S3A                                                                       ,7A                                                                                                                                                                                                                                                           �2A                        �         89A                       �         C9A                                  �1A                                   3A     !                             S3A     "                                     $                             �7A     %                                    &                            3A     '                            ��@     (                                    )                            ��@     *                                    +                            �@     ,                             �2A                                          .                                     !                  �         89A     0                  	�         C9A                                  �1A     1                             3A     2                             S3A     3                             x8A     5                            x8A     6                             �2A     1                   �         89A                       �         C9A                    	              �1A     9               	              3A     :               	              S3A     ;               	             �3A     =               	             W5A     >               	              �2A     9               
    �         89A     @               
   �                 A               
   �         C9A     B               
   �         C9A                                 �1A     D                            �1A     C                            3A     E                            S3A     F                             \4A     H                            \4A     I                             �2A     C                             �1A     J                             3A     K                             S3A     L                             �5A     N                            �2A     J                   �         89A                       �         89A                                  �1A     Q                             3A     R                             S3A     S                             �9A     U                     
       �3A     V                     
       }5A     W                            �2A     Q                   �         89A     Y                  �         C9A                                         [                                    \                                                         �                 ^                                    _                                    `                                                        �                 b                  �                 a                  �                 d                  �                 e                  �                                     �                 g                  �                 f                  �                 i                  �                 j                  �                                     �                 l                  �                 k                   �                 n                  �                 o                  �                 p                  �                 q                  �                                     �                 r                   �                 t                  �                 s                   �                 v                  �                 w                  �         N9A     x                  �                 y                  �                 z                  �                                     �                 |                  �                 }                  �                 ~                  �                                    �         ��@     �                  �                 �                  �                                     �                 �                  �                 �                   �                 �                  �                 �                  �                 �                  �                 �                  �                 �                  �                 �                  �                 �                  �                 �                  �                 �                  	�                                     �                 �                  �                 �                   �                 �                  �                 �                  �                 �                  �                 �                  �                                        ����                                                  �                                    �                                    �                                    �                                    �                  �                 �                                    �                            ��@     �                     
               �                     
       h�@     �                  	   
       ��@     �                  
   
               �                     
               �                     
               �                     ����                                                 �                            ��@     �                            ��@     �                                    �                                    �                                    �                                    �                                    �                     ����                                   
       ��@     �                     
       ��@     �                             f�@     �                             f�@     �                            f�@     �                            f�@     �                            f�@     �                            f�@     �                            f�@     �                            f�@     �                     
       ]�@     �                            ��@     �                                    �                                    �                            ��@     �                                    �                            g�@     �                  	          ��@     �                  
                  �                     ����                                                 �                            ��@     �                            ��@     �                                    �                                    �                                    �                                    �                                    �                     ����                               
                  �                  	                  �                                    �                                    �                      
       ��@     �                     
       ��@     �                             f�@     �                             f�@     �                            f�@     �                            f�@     �                            f�@     �                            f�@     �                            f�@     �                            f�@     �                     
       ]�@     �                  �  
       2�@     �                     
               �                                    �                            ��@     �                                    �                            g�@     �                  	          ��@     �                  
                  �                     ����                                                 �                            ��@     �                            ��@     �                                    �                                    �                                    �                                    �                                    �                     ����                                                 �                  
                  �                  	                  �                                    �                                    �                      
       ��@     �                     
       ��@     �                             ��@     �                             ��@     �                            ��@     �                            ��@     �                            ��@     �                            ��@     �                            ��@     �                            ��@     �                            ��@     �                            ��@     �                            ��@     �                            ��@     �                  �          7�@                       �  
       ]�@                      �         	�@                      �         ]�@                      	�         ]�@                      
�         ]�@                      �         ]�@                      �         ]�@                      �         ]�@                      �         [�@     	                 �                 �                  �  
                                �  
                                �  
               �                                                               ��@     �                                                               g�@                                ��@                                                                                                                                                                                                                                           ����                                 �         ��@                       �         A�@                        �         A�@                       �         A�@                       �         ��@                       �         A�@                       �         A�@                        �         A�@     !                  �         A�@     "                  �         A�@     #                  �         A�@     $                  �         A�@     %                  �         A�@     &                  �         A�@     '                  �         A�@     (                  �         A�@     )                  �         A�@     *                  �         A�@     +                  �         ��@     ,                  �         A�@     -                  �         A�@     .                  �         A�@     /                  �         A�@     0                  �         A�@     1                  �         A�@     2                  �         A�@     3                  �         A�@     4                  �         A�@     5                  �         A�@     6                  �         A�@                                          8                                   9                                   :                                   ;                                                   !    �         ��@     =              !   �         ��@     <              "    �                 ?              "   �                 @              "   �                                 #       
       ��@     B              #      
       ��@     A              #              f�@     D              #              f�@     E              #             f�@     F              #             f�@     G              #             f�@     H              #             f�@     I              #             f�@     J              #             f�@     K              #             f�@     L              #             f�@     M              #             f�@     N              #             f�@     C              #              ]�@     P              #             H�@     Q              #             ]�@     R              #             j�@     C              #   	�          ]�@     T              #   	�  
       ]�@     U              #   
   
       ��@     V              #   
   
       ]�@     C              #                     X              #             ��@     C              #                     Z              #                     [              #             g�@     \              #             ��@     ]              #                     ^              #      ����                            #                     `              #                     a              #                     b              #                     c              #                     d              #                     C              $    �                 f              $   �                 e                 �                 h                 �                 i                 �                                 %              ��@     k              %             ��@     j              %              f�@     m              %              f�@     n              %             f�@     o              %             f�@     p              %             f�@     q              %             f�@     r              %             f�@     s              %             f�@     t              %             f�@     u              %             f�@     v              %             f�@     w              %             f�@     l              %             H�@     y              %   �  
       _�@     z              %             ]�@     {              %             ]�@     |              %   �  
       ��@     }              %             ]�@     ~              %             ]�@                   %   �  
       ��@     �              %             ]�@     �              %             ]�@     l              %   	                  �              %   	          ��@     l              %   
                  �              %             g�@     �              %             ��@     �              %                     �              %                     �              %                     �              %                     �              %                     �              %                     �              %      ����    ��@                     %                     �              %                     �              %                     �              %                     �              %                     �              %                     �              %                     �              %   
                  l              &       
       ��@     �              &      
       ��@     �              &              f�@     �              &              f�@     �              &             f�@     �              &             f�@     �              &             f�@     �              &             f�@     �              &             f�@     �              &             f�@     �              &      
       ]�@     �              &   �         ��@     �              &   �         ��@     �              &             I�@     �              &                     �              &             ��@     �              &                     �              &             g�@     �              &   	          ��@     �              &   
                  �              &                     �              &                     �              &      ����                            &                     �              &             ��@     �              &             ��@     �              &                     �              &                     �              &      ����                            &                     �              &                     �              &                     �              &   
                  �              &   	                  �              &                     �              &                     �                      
       ��@     �                     
       ��@     �                             f�@     �                             f�@     �                            f�@     �                            f�@     �                            f�@     �                            f�@     �                            f�@     �                            f�@     �                            ]�@     �                            ]�@     �                            �@     �                                    �                            ��@     �                                    �                  	          g�@     �                  
                  �                            ��@     �                     ����                                                  �                            ��@     �                                    �                            ��@     �                                    �                                    �                                    �                     ����                                                  �                                    �                  
                  �                  	                  �                                    �              '       
       ��@     �              '      
       ��@     �              '              f�@     �              '              f�@     �              '             f�@     �              '             f�@     �              '             f�@     �              '             f�@     �              '             f�@     �              '             f�@     �              '             ]�@     �              '             ]�@     �              '             k�@     �              '                     �              '             ��@     �              '                     �              '   	          g�@     �              '   
                  �              '             ��@     �              '                     �              '      ����                            '                     �              '                     �              '                     �              '   
                  �              '   	                  �              '                     �              (       
       ��@     �              (              f�@     �              (             ]�@     �              (             ]�@     �              (   �         ��@     �              (                     �              (             ��@     �              (                     �              (                     �              (             g�@                    (                                   (   	                                (   
          ��@                   (      ����                            (                                   (   
                                (   	                                (                                   (                     	              (                     �              )    �                               )   �                 
              )   �                               )   �                               )   �                                 *       
       ��@                   *      
       ��@                   *              f�@                   *              f�@                   *             f�@                   *             f�@                   *             f�@                   *             f�@                   *             f�@                   *             f�@                   *             ]�@                   *             ]�@                   *             7�@                   *                                   *             ��@                   *                                   *   	          g�@                    *   
                  !              *             ��@     "              *                     #              *                     $              *      ����    ��@                     *                     &              *                     '              *                     (              *                     )              *   
                  *              *   	                  +              *                                   +       
       ��@     -              +      
       ��@     ,              +              f�@     /              +              f�@     0              +             f�@     1              +             f�@     2              +             f�@     3              +             f�@     4              +             f�@     5              +             f�@     .              +             ]�@     7              +             ]�@     8              +             7�@     .              +                     :              +             ��@     .              +                     <              +   	          g�@     =              +   
                  >              +             ��@     ?              +                     @              +                     A              +      ����                            +                     C              +                     D              +                     E              +                     F              +   
                  G              +   	                  H              +                     .              ,    �  
       ��@     J              ,   �  
       ��@     I              ,    �         f�@     L              ,   �         f�@     K              ,   �  
       ]�@     N              ,   �         `�@     O              ,   �                 P              ,   �                 O              ,   �                 R              ,   �         ��@     K              ,   �                 T              ,   �         g�@     U              ,   �                 V              ,   �         ��@     W              ,   	                  X              ,   
                                  -       
       ��@     Z              -      
       ��@     Y              -              ��@     \              -              f�@     ]              -             f�@     ^              -             f�@     _              -             ��@     `              -             f�@     a              -             f�@     b              -             f�@     c              -             ��@     d              -             f�@     e              -             f�@     f              -             f�@     [              -    �         ]�@     h              -   �         2�@     i              -   �         2�@     j              -   �         ��@     h              -                     l              -             ��@     [              -   	          g�@     n              -   
   
       ��@     o              -      
               p              -      
               q              -      
               r              -      
               s              -      
               t              -      
               u              -      
               v              -                     w              -      ����    ��@                     .       
       ��@     y              .      
       ��@     x              .                      {              .              ��@     |              .              f�@     }              .             f�@     ~              .             f�@                   .             f�@     �              .             f�@     �              .             ��@     �              .             f�@     �              .             f�@     �              .             f�@     �              .             f�@     �              .             f�@     {              .    �         ]�@     �              .   �         ��@     �              .   �                 �              .   �         ��@     �              .                     �              .             ��@     {              .   	          g�@     �              .   
          ��@     �              .                     �              .                     �              .                     �              .                     �              .      ����    ��@                     .                     �              .                     �              .                     �              .                     �              .                     �              .   
                  �              .   	                  {              /    �                 �              /   �                 �              0    �                 �              0   �                 �              0   �                 �              0   �                 �              0   �                                 1       
       ��@     �              1      
       ��@     �              1              ��@     �              1              f�@     �              1             f�@     �              1             f�@     �              1             f�@     �              1             f�@     �              1             ��@     �              1             f�@     �              1             ]�@     �              1             �@     �              1             ]�@     �              1             �@     �              1             ]�@     �              1             �@     �              1      
       ��@     �              1      
               �              1      
       g�@     �              1   	   
               �              1   
   
               �              1      
               �              1      
       ��@     �              1      
               �              1      
               �              1                     �              1      ����    ��@                     2       
       ��@     �              2              f�@     �              2              f�@     �              2             f�@     �              2             f�@     �              2             f�@     �              2             f�@     �              2             ]�@     �              2             ]�@     �              2   �         ]�@     �              2   �          �@     �              2                     �              2             ��@     �              2   �                 �              2   �         g�@     �              2   	�                 �              2   
�                 �              2   �         +�@     �              2   �                                 2                     �              2                     �              2   
                  �              2   	                  �              2                     �              2                     �              3       
       ��@     �              3      
       ��@     �              3              f�@     �              3              f�@     �              3             f�@     �              3             f�@     �              3             f�@     �              3             f�@     �              3             f�@     �              3             f�@     �              3      
       ]�@     �              3      
       ]�@     �              3   �         ��@     �              3             ]�@     �              3   �         ��@     �              3             I�@     �              3                     �              3             ��@     �              3                     �              3   	          g�@     �              3   
          ��@     �              3                     �              3      ����                            3                     �              3             ��@     �              3             ��@     �              3                     �              3                     �              3                     �              3                     �              3                     �              3      ����                            3                     �              3                     �              3   
                  �              3   	                  �              3                     �              4       ����            �              4                      �              4                     �              4             g�@     �              4                                    4                                   4                                   4                                   4                                   4                                   4   	                                4   
          A�@                   4      ����                            4                     	              4             ��@     �              5       ����                            5      $       ��@     
              5       d       ��@                   5       
                             5       
                             5       ����    ��@                     3       
       ��@                   3       �       &�@                   3       �       ��@                   6    �         Q�@                   6   �         I�@                   6   �         I�@                   6   �         I�@                        �         A�@                       �         A�@                       �         A�@                       �         A�@                       �         A�@                       �         A�@                       �         A�@                       �         A�@                        �  
                                 �  
               !                 �  
       =�@                     7                      #              7   �                 "              8                      %              8   �                 $              9                      '              9                     &              :    �                 )              :   �         g�@     *              :   �                 +              :   �  
       ��@     ,              :   �  
                               ;    �                 .              ;   �                 /              ;   �                 -              <                      1              <                     2              <                     3              <                     4              <                     5              <                     0              =                      7              =                     8              =                     9              =                     :              =                     ;              =                     6              >       
               =              >   �  
               <              ?       
               ?              ?   �  
               >              @       
               A              @   �  
               @              A       
               C              A   �  
               B              B       
               E              B   �  
               D              C       
               G              C   �  
               F              D       ����                            E       ����                            F    �                 K              F   �                 L              F   �                 M              F   �                 N              F   �                 O              F   �                 J              G    �                 Q              G   �                 R              G   �                 S              G   �                 P              H    �  ����                            I    �                 V              I   �                 W              I   �                 X              I   �                 U              J    �                 Z              J   �                 [              J   �                 \              J   �                 Y              K    �  ����                            L    �                 _              L   �                 `              L   �                 a              L   �                 b              L   �                 c              L   �                 ^              M    �                 e              M                     d              N       ����                            O       ����                            P       ����                            Q       ����                            R       ����                            S       ����                            T       ����                            U       ����                            V       ����                            W       ����                            X       ����                            Y       ����                            Z       ����                            [       ����                            \       ����                            ]       ����                            ^    �  ����                            _       ����                            `       
               y              `                     z              `                     {              `                     x                    ����                                  ����                            a       ����                            b       ����                            c       ����                            d    �                 �              d   �                 �              e       ����                            f                      �              f                     �              g       ����                            h       ����                            i       ����                            j       ����                            k       ����                            l       ����                            m       ����                            n       ����                            o       ����                            p    �  ����                            q    �  ����                            r       ����                            s       ����                            t       ����                            u       ����                            v    �                 �              v   �                 �              v   �                 �              v   �                 �              w    �                 �              w   �                 �              w   �                 �              x                      �              x                     �              y    �                 �              y   �                 �              y   �                 �              y   �                 �              z    �                 �              z   �                 �              z   �                 �              z   �                 �              {    �                 �              {   �                 �              {   �                 �              {   �                 �              |    �                 �              |   �                 �              |   �                 �              |   �                 �              }    �                 �              }   �                 �              }   �                 �              }   �                 �              ~    �                 �              ~   �                 �              ~   �                 �              ~   �                 �                     ����                            �       ����                            �       ����                            �       ����                            �       ����                            �       ����                            �       ����                            �       ����                            �       ����                            �    �                 �              �   �                 �              �   �                 �              �   �                 �              �    �                 �              �   �                 �              �   �                 �              �   �                 �                      ӐB     ؐB     ݐB     �B     �B     �B     �B     ��B     ��B      �B     �B     
�B     �B     �B     �B     �B     #�B     (�B     -�B     2�B     7�B     <�B     A�B     F�B     K�B     P�B     U�B     Z�B     _�B     d�B     i�B     �aB     n�B     s�B     x�B     }�B     ��B     ��B     ��B     ��B     ��B     ��B     ��B     ��B     ��B     ��B     ��B     ��B     ��B     ÑB     ȑB     ͑B     ґB     בB     ܑB     �B     �B     �B     �B     ��B     ��B     ��B     �B     	�B     �B     �B     �B     �B     "�B     '�B     FaB     ,�B     1�B     6�B     ;�B     @�B     E�B     J�B     O�B     T�B     O�B     Y�B     ^�B     c�B     h�B     m�B     r�B     w�B     |�B     ��B     ��B     ��B     ��B     ��B     ��B     ��B     ��B     ��B     ��B     ��B     ��B     ��B     B     ǒB     ̒B     ђB     ֒B     ےB     ��B     �B     �B     �B     ��B     ��B     ��B     �B     �B     �B     �B     �B     �B     !�B     &�B     +�B     0�B     5�B     :�B     ?�B     D�B     I�B     N�B     S�B     X�B     ]�B     b�B     g�B     l�B     q�B                                                 	   ����   ����          |�B           D�             h�B                             @8e     w                       B�B                             T�B                             n�B                             y�B                             ��B                             ��B                             ��B                             ��B                             B                             ̗B                             ӗB                            �B                             ��B                             �B                             �B                             '�B                            4�B                            �RB                             @�B                             �RB                             �RB                             P�B                             i�B                            v�B                            ��B                             ��B                             ǓB                             ��B                             ٓB                             ��B                             �B                             ��B                             ��B                             ��B                             ԘB                             �B                             �B                             "�B                             <�B                             V�B                             p�B                             ��B                             ��B                             ��B                             ��B                             ΙB                             ޙB                             �B                             �B                             �B                             �B                             0�B                             B�B                             M�B                            W�B                            i�B                            u�B                            ��B                            ��B                            ��B                            ��B                            ��B                            КB                            ߚB                            �B                            ��B                            	�B                            �B                            )�B                            8�B                            I�B                            [�B                            j�B                            x�B                            ��B                            ��B                            ��B                            ��B                            ɛB                            ؛B                            �B                            ��B                            �B                            �B                            �B                            -�B                            =�B                            L�B                            Y�B                            f�B                            x�B                            ��B                            ��B                            ��B                            ��B                            ��B                            ��B                            ̜B                            ؜B                            �B                            ��B                            �B                            �B                            &�B                            ;�B                            M�B                            d�B                            q�B                            ��B                            ��B                            ��B                            ��B                            ϝB                            �B                            ��B                            �B                            #�B                            8�B                            M�B                            @Ge     L                       SRB                             eRB                             pRB                             b�B                             l�B                             }RB                             y�B                            ��B                            ��B                            ��B                            ��B                            ��B                            ��B                            ɞB                            ҞB                            ܞB                            �B                            ��B                            �B                            �B                            �B                            *�B                            6�B                            A�B                            L�B                            X�B                            c�B                            o�B                            |�B                            ��B                            ��B                            ��B                            ��B                            ��B                            ǟB                            ԟB                            ݟB                            �B                            �B                            ��B                             �B                             �B                             �B                             -�B                             v�B                             9�B                             C�B                             O�B                             X�B                             c�B                             �RB                             m�B                             �RB                             �RB                             x�B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ȠB                            РB                             ۠B                            �B                            �B                            ��B                            �B                            �B                            �B                            %�B                            0�B                            ;�B                            F�B                            Q�B                            \�B                                ������������������������         -   =   �   �   �   �   �   �   �   �   �   �   �   n   y         �   �   �   �      c   m   g   f   0   	   -   =   �   �   �   �   8   7   6   5   4   3   2   1   t   �   q   �      ����������������������������            �   �   k   z   w   q   h   5   6   7   8   9   0   \      /      ]   [   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �       P   ]   _      8   H   N   4   9            #   $   &   4           Ye     �Re     �@     P 6                                            8�@     1                      8�@     2                      8�@     3                      8�@     4                      8�@     5                      8�@     6               Ye     �Se     ��@     P 6                                            �@     1                      �@     2                      �@     3                      �@     4                      �@     5                      �@     6               Ve     �Te     ��@     P @                              M_SFXVOL      i�@     s       ��                               M_MUSVOL      ��@     m       ��                                     �Ue     �Ue     Q�@     J�                                            ��@                     Ye      Ve     ��@     �                                            ��@                     Ye     `Ve     �@     < %                              M_ENDGAM      ע@     e        M_MESSG       �@     m        M_DETAIL      ל@     g        M_SCRNSZ      ,�@     s       ��                               M_MSENS       ~�@     m       ��                               M_SVOL         �@     s              @Xe     �We     ��@     0 ?                             M_JKILL       m�@     i        M_ROUGH       m�@     h        M_HURT        m�@     h        M_ULTRA       m�@     u        M_NMARE       m�@     n               Ye     �Xe     ߚ@     0 ?                              M_EPI1        K�@     k        M_EPI2        K�@     t        M_EPI3        K�@     i        M_EPI4        K�@     t                      @Ye     x�@     a @                              M_NGAME       
�@     n        M_OPTION      ��@     o        M_LOADG       �@     l        M_SAVEG       4�@     s        M_RDTHIS      ��@     r        M_QUITG       �@     q       ��B     ħB                     Gamma correction OFF      Gamma correction level 1  Gamma correction level 2  Gamma correction level 3  Gamma correction level 4    
                                                            ��     ��      hH��  ��hH��   ��      hH��  ��hH��    ��                                                                      
            �   2   ,  2                                                      NUKAGE3  NUKAGE1           FWATER4  FWATER1           SWATER4  SWATER1           LAVA4    LAVA1             BLOOD3   BLOOD1            RROCK08  RROCK05           SLIME04  SLIME01           SLIME08  SLIME05           SLIME12  SLIME09          BLODGR4  BLODGR1          SLADRIP3 SLADRIP1         BLODRIP4 BLODRIP1         FIREWALL FIREWALA         GSTFONT3 GSTFONT1         FIRELAVA FIRELAV3         FIREMAG3 FIREMAG1         FIREBLU2 FIREBLU1         ROCKRED3 ROCKRED1         BFALL4   BFALL1           SFALL4   SFALL1           WFALL4   WFALL1           DBRAIN4  DBRAIN1       ����                                                    SW1BRCOM SW2BRCOM  SW1BRN1  SW2BRN1   SW1BRN2  SW2BRN2   SW1BRNGN SW2BRNGN  SW1BROWN SW2BROWN  SW1COMM  SW2COMM   SW1COMP  SW2COMP   SW1DIRT  SW2DIRT   SW1EXIT  SW2EXIT   SW1GRAY  SW2GRAY   SW1GRAY1 SW2GRAY1  SW1METAL SW2METAL  SW1PIPE  SW2PIPE   SW1SLAD  SW2SLAD   SW1STARG SW2STARG  SW1STON1 SW2STON1  SW1STON2 SW2STON2  SW1STONE SW2STONE  SW1STRTN SW2STRTN  SW1BLUE  SW2BLUE   SW1CMT   SW2CMT    SW1GARG  SW2GARG   SW1GSTON SW2GSTON  SW1HOT   SW2HOT    SW1LION  SW2LION   SW1SATYR SW2SATYR  SW1SKIN  SW2SKIN   SW1VINE  SW2VINE   SW1WOOD  SW2WOOD   SW1PANEL SW2PANEL  SW1ROCK  SW2ROCK   SW1MET2  SW2MET2   SW1WDMET SW2WDMET  SW1BRIK  SW2BRIK   SW1MOD1  SW2MOD1   SW1ZIM   SW2ZIM    SW1STON6 SW2STON6  SW1TEK   SW2TEK    SW1MARB  SW2MARB   SW1SKULL SW2SKULL                                                                                                                                                                                                          @  ����@  ����@  @  ����@  @  ����@  @  @  ����@  @  @  ����������������@  ��������@  @  @  @  ����@  ����@  @  ��������@  @  ����������������@  @  @  @  ����@  @  ����@                                 none                    ��������        ����                    pistol      @           ��������        ����                    shotgn      @           ��������        ����                    sgcock      @           ��������        ����                    dshtgn      @           ��������        ����                    dbopn       @           ��������        ����                    dbcls       @           ��������        ����                    dbload      @           ��������        ����                    plasma      @           ��������        ����                    bfg         @           ��������        ����                    sawup       @           ��������        ����                    sawidl      v           ��������        ����                    sawful      @           ��������        ����                    sawhit      @           ��������        ����                    rlaunc      @           ��������        ����                    rxplod      F           ��������        ����                    firsht      F           ��������        ����                    firxpl      F           ��������        ����                    pstart      d           ��������        ����                    pstop       d           ��������        ����                    doropn      d           ��������        ����                    dorcls      d           ��������        ����                    stnmov      w           ��������        ����                    swtchn      N           ��������        ����                    swtchx      N           ��������        ����                    plpain      `           ��������        ����                    dmpain      `           ��������        ����                    popain      `           ��������        ����                    vipain      `           ��������        ����                    mnpain      `           ��������        ����                    pepain      `           ��������        ����                    slop        N           ��������        ����                    itemup      N           ��������        ����                    wpnup       N           ��������        ����                    oof         `           ��������        ����                    telept                  ��������        ����                    posit1      b           ��������        ����                    posit2      b           ��������        ����                    posit3      b           ��������        ����                    bgsit1      b           ��������        ����                    bgsit2      b           ��������        ����                    sgtsit      b           ��������        ����                    cacsit      b           ��������        ����                    brssit      ^           ��������        ����                    cybsit      \           ��������        ����                    spisit      Z           ��������        ����                    bspsit      Z           ��������        ����                    kntsit      Z           ��������        ����                    vilsit      Z           ��������        ����                    mansit      Z           ��������        ����                    pesit       Z           ��������        ����                    sklatk      F           ��������        ����                    sgtatk      F           ��������        ����                    skepch      F           ��������        ����                    vilatk      F           ��������        ����                    claw        F           ��������        ����                    skeswg      F           ��������        ����                    pldeth                  ��������        ����                    pdiehi                  ��������        ����                    podth1      F           ��������        ����                    podth2      F           ��������        ����                    podth3      F           ��������        ����                    bgdth1      F           ��������        ����                    bgdth2      F           ��������        ����                    sgtdth      F           ��������        ����                    cacdth      F           ��������        ����                    skldth      F           ��������        ����                    brsdth                  ��������        ����                    cybdth                  ��������        ����                    spidth                  ��������        ����                    bspdth                  ��������        ����                    vildth                  ��������        ����                    kntdth                  ��������        ����                    pedth                   ��������        ����                    skedth                  ��������        ����                    posact      x           ��������        ����                    bgact       x           ��������        ����                    dmact       x           ��������        ����                    bspact      d           ��������        ����                    bspwlk      d           ��������        ����                    vilact      d           ��������        ����                    noway       N           ��������        ����                    barexp      <           ��������        ����                    punch       @           ��������        ����                    hoof        F           ��������        ����                    metal       F           ��������        ����                    chgun       @   �ce     �               ����                    tink        <           ��������        ����                    bdopn       d           ��������        ����                    bdcls       d           ��������        ����                    itmbk       d           ��������        ����                    flame                   ��������        ����                    flamst                  ��������        ����                    getpow      <           ��������        ����                    bospit      F           ��������        ����                    boscub      F           ��������        ����                    bossit      F           ��������        ����                    bospn       F           ��������        ����                    bosdth      F           ��������        ����                    manatk      F           ��������        ����                    mandth      F           ��������        ����                    sssit       F           ��������        ����                    ssdth       F           ��������        ����                    keenpn      F           ��������        ����                    keendt      F           ��������        ����                    skeact      F           ��������        ����                    skesit      F           ��������        ����                    skeatk      F           ��������        ����                    radio       <           ��������        ����                                            1�B                             6�B                             ;�B                             @�B                             E�B                             J�B                             O�B                             T�B                             Y�B                             ^�B                             c�B                             h�B                             m�B                             r�B                             w�B                             |�B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             }YB                             ��B                             ��B                             �B                             �B                             �B                             �B                             �B                             CTB                             "�B                             )�B                             0�B                             6�B                             =�B                             D�B                             K�B                             R�B                             Y�B                             `�B                             f�B                             m�B                             t�B                             {�B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             ��B                             �  ��������                   idmypos                                                                                        idclev                                                                                        idchoppers                      
                                                               idbeholdv                       	                                       idbeholds                       	                                       idbeholdi                       	                                       idbeholdr                       	                                       idbeholda                       	                                       idbeholdl                       	                                       idbehold                                                                       idclip                                                                                         idspispopd                      
                                                               idfa                                                                                           idkfa                                                                                          iddqd                                                                                          idmus                                                                 ����         �C               h   �                                                                 (   �                                                                 �   `                                                                 h   P                                                                 x                                                                     (                                                                                    �   �                                                               �   �                                                               �   �                                                               �   �                                                               �   �                                                               �   �                                                               �   �                                                               �   �                                                               �   �                                                                                        �   h                                                                 �   �                                                                 p   �                                                                 H   p                                                                 X   `                                                                 @   0                                                                 �   (                                                                 �                                                                    P                                                                    @                                                          g)B     Q)B     )B        
      @   GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o ,             �@     -                       ,           ]@                            ,    �       ^@     �                          /l                           ��                       ,    �       [&@     d                           ֡                       ,    �       �&@     �                      ,    5�       �*@     q                      ,    ��       �/@     �                      ,    N[      �C@     *                      ,    �_      �D@     �                      ,    w�      dH@     �
                      ,    ��      JS@     J                      ,    ��      �W@     Q"                      ,    �t      �y@     �                      ,    >�      �~@     �                          �                      ,    73              #                       ,    �5      p�@                            ,    8      q�@     �                       ,    v<              �                      ,    �g      ,�@     9                      ,    �v      e�@                           ,    ׆      }�@     X                       ,    �              �                      ,    M�      Ս@     �                       ,    ��      [�@     =                       ,    ��      ��@     �                       ,    ]�      8�@     8                      ,    �      p�@     J                      ,    �      ��@     L                       ,    G�      �@     �                      ,    u=      ��@     �                      ,    sQ      ��@     G                       ,    lR      �@     B                      ,    0�      )�@     �                      ,    ��      ��@     �                      ,    �s      ��@     �                      ,    (�      �@                           ,    �!      0�@     �                      ,    *k      ��@     a                      ,    �      5A     `
                      ,    �-      �A     B                      ,    ތ      �*A     �                      ,    e�      �.A     �                      ,    �=      t:A     �                      ,    ��      .QA                           ,    �	      9^A     #                      ,    `	      \bA                           ,    ��	      joA                           ,    i
      �tA     �                      ,    c
      vA     �                       ,    H�
      wA     ~                      ,    ��
      �{A                           ,    t@      ��A     U                      ,    ��      ��A     =                      ,    G�      2�A     J	                      ,    �<      |�A                           ,    ��      ��A     �                      ,    �      +�A                            ,    _      6�A     �                      ,    _[      ��A     l                          Aa                      ,    �e      ]�A     E                       ,    :�      ��A     �                      ,    	�      0�A     �                      ,    E@      ��A     �                      ,    d�      ��A     )                       ,    q�      ��A     s                      ,    �      hB     �                      ,    R&      \B                           ,    �,      ^B     '                       ,    t0      �B     k                       ,    �4      �B                            ,    �F      �#B     /                      ,    �P      )B     �                       ,    V      �)B     �                       ,    |_      g*B     �                      ,    um      �.B                            <    �n      /B     
      @                            ,    I�      1B     u                       ,    �      �1B     E                      �    ��      �>B     �      �DB     2       �DB     �       vEB            �EB     -       �EB     -       �EB             FB     �       �FB     "       �FB     "       �FB     �       �GB     -                      ,    �      �HB     �                       ,    f�      �IB     �                                              S#  �  �*                      �)  �9   ,	  ^&  �  �1  @�   Q  �    �   	-   62  #	-     &	-   �5  )	-    �@  ,	-   (.  -	-   0*  2�   8;:  5�   < �   1  int �K 8"N   �  K�   �   �  L�   �  M�   e2    �0  }  �  �   q  O  �   	`R (�   �@     -       ��  
�  (�          
s  (O  A   =   �@     �  �@     �  �  U	�JB      @     �  	@     	   �  �  #     �  �  %�  �  ! �    �   S#  �C  �*  ]@            �  �  ,	  e2    �  �0  }  int ^&  F   J�   D   �C  
D  ���� �C  Ni   �C  	�   	T�e     �C  	�   	P�e     	�C  +]@            � 5i   �  S#  �[  �*  ^@     �      �  u  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �  	"|  *y  	��  +y  	I�  ,y  	�a  -y  
K   "  ��  WH  �~  �O  �m  ��   �  ��  ��  	 
K   	V  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  	(  
K   	/�  ��   [r  �4 #�  �   �X  	5b  
K   	:�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  	K�  
�   	P=  =_  ��   R�  N�  ��  ��   �p  	W
  
K   
3p  ��   ({  ��  ğ   F]  
8I  
K   
Y�  ��   �c  |  ��  l  ��  �   
K   
k  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  
{�  
K   
�E  &�   �  º  GY  �f  ��   v�  
�  
K   
��  GQ   ϼ  �  �_  X  &�  �b   
K   !�  �p   �  ��  S�  ��   �F  '�  *	  *� ,�   "G  C	�   (G  C�   �]  C�   :G  C�    �U  D�  H#	r  � '
r   �^  (1    .�  )	�   (o�  -1   0i�  .	�   8��  /
�  < �   �  =    �   �  =    �  0  	p�  L�  �  	t�  M�  	K�  N�  	x�  O�  	��  P�  	��  Q�  	r�  R�  �    =    	�  S�  	�u  T�  		�  U�  	h�  V�  t�   �   8  D  Z  =   �' I  	��  1Z  	]  4w  D  D  �  =   � }  	Zy  8�  �  �  =   =   � �  	��  ;�  Ʃ  QK   �  �  �  =     �  	�  W�  �p  #       S�  $  $  /  R    T}  %;  A  Q  R   R    '	  acv )�  ��  *  ��  +/   �y -Q  �Y  6  ��  :�  s�  <�   �H  =�  xz  >�   �  x @�  �   �  =    B  �  =    4    =    
�	U  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x �  
K   �  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �a  
K   �E%  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�  (x	�%  �u z�   � {	�   s |	�   � ~  N�  E%  ��  �	�   ��  �	�     J]  �R%  �%  �%  =   � �^  ��%  �   �%    �  ��%  !K   �N)  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  &  \	�*  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /[)  �*  �*  =   � ��  1�*  �]  ���,  `e ��   x �8  y �8  z �8   ��  ��,  (cN  ��,  0Mp ��  8�u ��  <� ��   @�H  ��,  Hr�  ��,  P��  ��,  X��  �8  `m�  �8  d��  �8  h  �8  l3F  �8  p8F  �8  t=F  �8  x��  ��   |*� �N)  �y� ��,  �s ��   ��� ��,  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  �,  ���  �   ���  	�   ��R  �.  �f�  �   �I}  U  ���  �,  � �*  Gx  ��,  >} ��2   �}  �B  �|  �B  
 �,  �*  �%  "d  HN�.  mo PN1   ��  Q�8  cmd R�8  �  W8  (_  Y8   #_  [8  $bob ]8  (�  a�   ,�[  b�   0sb  d�   4d]  g�8  8�W  h�8  P��  iy  h�� lT1  l�N  m  |E�  p  ��W  r9  �~�  sT1  �*� tT1  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �N1  �#�R  ��    #��  ��   #�  ��   #h  �9  #I�  �y  @ �,  �z �*  	��  ��   	�\  �y  	�  �/  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  ��  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   (	�/  ��  B      B  Vd  !B  �  "B  �� #�/   �   �/  =    � %�/  C	$0  x E8   y F8   �{ H0  (T	h0  `e V�   x W8  y X8  z Y8    	�  [00  �a	N1  = c8   F�  d8  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  oN1  ��  r
T1   iK  uh0  0��  x
�   XS�  {N1  `��  ~R   h��  ��   pu| �$2  x �.  �   d1  =    �}  X�$2  v1 ��2   v2 ��2  dx �8  dy �8  �  �B  �k �B  tag �B  �W  ��  �o ��2  $��  ��2  4SX  ��2  8d�  ��2  @��  �
�   H��  �R   P *2  d1  �z �t0  �	�2  2�  �8   ]  �8  �h  �B  �N  �B  
�K  �B  >} ��2   02  �}  �<2  
K   ��2  ��   �  o�  ��   ��  ��2  $0  8  �2  =    �u  �d1  �z ��,  8�	w3  v1 ��2   v2 ��2  82  �8  Mp ��  [�  �w3   �  �}3   SX  ��2  (d�  ��2  0 �2  �2  A{ �3  4	�3  $x 8   $y 	8  $dx 
8  $dy 8  �o �3  )�  �  0 8  �3  =   =    (} �3  �  *�  %v  @2�4  @�  4�4   $x1 5�   $x2 6�   .]  88  5]  98  �� :8  ��  =�   �  @8   ��  C8  $�n  G�4  (9x  H�4  0�^  I�4  8 �3  B  >�  K4  %�h  PR�5  s�  U�5   �H  V�5  $x1 X�   $x2 Y�   $gx \8  $gy ]8  $gz `8   $gzt a8  $�x  d8  (� f8  ,~�  i8  0t  k8  4.� l�   8�  p�5  @	�  r�   H �4  4  �h  t�4  �	6  �c  �y   �O  �6  �x  �
 6   B   6  =    �  06  =    I�  ��5  �	d6  �  ��    �  �d6   06  �  �=6  &��	!7    �8   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  $top �	!7  '��  �	�  U'��  �	�  V'� �	!7  W'�  �	�  � �  27  =   ? ��  �w6  	�7  ~�  E   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %?7  �7  �7  =    	S�  '�7  
K   7�7  {�   U�  ~�   >	8  �� @�,   s A
�   sx B8  sy C8   Nz E�7   	�8  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4(8  
K   1�8  ��   ��  ��   �y  9�8  �   �8  =    y  9  =    y  9  =    8  -9  =    hy ��,  (�	�9  in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
T1  �a  �
�   $ ��  �99  ��	B:  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  �B:  ( �9  R:  =    ޴  ��9  	.L  &j:  8  	׮  )j:  	�  +j:  	�  ,j:  	�Q  .�5  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�:  �   	��  8�:  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F*;  j6  	��  H�   	��  I�2  	��  K�   	a� L�4  	w�  N�   	P{ O�2  	��  Q�   	��  R�;  �2  	��  T�   	�� U�;  �3  	�}  W�   	u| X}3  	M�  Z�   	P�  [w3  	��  a8  	��  b8  	�  c8  	�p  e�  	�T  f <  -9  	�a  j�  �   C<  =   � 	ը  l2<  �  `<  =   @ 	�p  mO<  	 �  p8  	p|  q�  	$Y  v�   	�K  y�   	g  {�<  27  	d�  |�<  	��   8  		�  !8  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +8  	`�  ,8  	A�  -8  	��  /�   	��  1�   	P�  2�   �5  `=  =   =   / 	��  EJ=  �5  |=  =   / 	Ԁ  Fl=  �5  �=  =   =    	7� G�=  	�R  I�   	��  J�5  	��  U�   (	P�  \�=  �=  	��  ]�=  	L�  ^�=  	ߵ  _�=  	�  a�=  	@�  �4  	[�  w3  	 �  }3  	SX  �2  	d�  �2  	��  �   	_�   �   	��  "y  	��  %y  	'�  &y  	�]  (y  �4  �>  =   � 	�P  *�>  	ӯ  +�>  �4  	|  -�>  �5  	��  .�>  	��  /�>  �>  ?  �   �    	��  �4  �   �>  	qY  "?  	�  #?  B  D?  =   ? 	��  %3?  	��  &3?  8  l?  =   � 	@Y  (\?  8  �?  =   ? 	V�  )x?  �5  �?  =    	�h  �?  	�  �?  �5  	�  �5  	�f  !3?  	r�  "3?  	��  %�4  	��  &�4  	׆  '8  	��  (8  	�  *8  	��  +8  	�   �5  	��   �   	�_   �   	�_   �   	b   8  	t   8  	j�   "�  	�   :�   	��   ;�   	��   <�   	�W   >�5  	hn   @8  	U~   A8  	�   B8  	 �   C8  	%�   F�  	�u   H�  	z   I�  	ʓ  !C�  U  #A  =    	��  !bA  �   ?A  =    	��  !c/A  	0K  !d�   	?�  !e�   !�	�A  x !�8   y !�8  dx !�8  dy !�8   ��  !�cA  !��A  �p !�
N1  ��  !�
}3   !�	�A  {q !�8   ��  !�y  d !�	�A   t�  !��A  �A  B  =   � 	r !�B  	�T  !�,B  �A  	l�  !�8  	�  !�8  	?k  !�8  	�d  !�8  	2~ !��A  	��  !�y  	��  !�8  	k�  !�8  	Z�  !�}3  }3  �B  =    	�v  !��B  	�v  !��   	"�  !�N1  �  !�  �U  !�4  ��  !�4  t�  !�   �  !	�   .Y  !
8  7Y  !8  �h  !:C  N1  *� !T1  <i  !T1  	G  "y  	��  "�   �   �C  =    
K   "��C  )top  �G  �  �]  "��C   "�	�C  ��  "�}3   ��  "��C  O{  "�
�   ��  "�
�   iK  "��C   h0  ��  "��C   D  D  =    	��  "�D  !K   "OD  )up  �  �F  �S   FT  "
(D  !K   "�D  ��   �x  H�  ��  �H   ��  "\D  H"	JE  `e "�   >} "�2  L� "8   $low "8  $+� " 8  (�Z "!
�   ,r� ""
�   0�f  "#OD  4�f  "$OD  8��  "%y  <$tag "&
�   @*� "'�D  D �w ")�D  gE  gE  =    JE  �  "2WE  !K   "��E  ��   �s  z�  ��  �T  ܭ   gY  "�zE  H"�	RF  `e "��   *� "��E  >} "��2   �W  "�8  (�}  "�8  ,L� "�8  0��  "�y  4��  "�
�   8$tag "�
�   <��  "�
�   @  w "��E  oF  oF  =    RF  j�  "_F  =� #�F  ��  #.�F  ^�  #2PG   }�  #7�  �� #;K    #	�F  r� # 	G   .� #$G  O� #)>G   *G  G  �    �F  �F  G  G   G  *1   >G  G  K   R   1     G  ��  #,�F  DG  oS  $'bG  dS  ($)�G  � $+
�   � $,G  @�  $-
�   >z $.
�   �  $/R   �H  $3�G    VG  	�� $7�G  	�� $8K   	<]  %�   	��  %�   	h  %�   	��  %�   	�  %�   	�j  %�   	��  %�   	v  %�   	R  %�   	��  %�   	�o  % �   	�U  %"�   	�n  %#�   	�  %$�   	��  %%�   	�  %&�   	��  %'�   	u  %(�   	_b  %)�   	N  %*�   	�  %-�   	��  %.�   	0h  %/�   	�g  %0�   	��  %1�   	^�  %2�   	�a  %3�   	>�  %4�   	��  %5�   	O  %7�   	��  %8�   	Ϊ  %:�   	��  %;�/  	ӄ  %=�   	r�  %>�   	~�  %?�   	��  %@�   	��  %A�   	��  %B�   	��  %C�   	��  %D�   	�T  %F�   		�  %G�   	^�  %H�   	��  %I�   	��  %J�   	�  %K�   	[n  %L�   	��  %M�   	-�  %O�   	��  %P�   	��  %Q�   	J�  %R�   	Ei  %T�   	��  %U�   	��  %V�   	A�  %W�   	��  %X�   	��  %Y�   	��  %Z�   	 t  %[�   	��  %\�   	!�  %]�   	oa  %^�   	/z  %_�   	��  %c�   	1P  %d�   	�  %e�   	Ʒ  %f�   	�T  %g�   	�o  %h�   	�b  %i�   	~�  %j�   	��  %k�   	�S  %m�   	��  %n�   	U  %o�   	Dl  %p�   	��  %q�   	��  %r�   	�p  %s�   	"�  %t�   	�  %u�   	�K  %v�   	��  %w�   	�  %y�   	tW  %z�   	'�  %{�   	��  %}�   	��  %~�   	�P  %�   	#L  %��   	gz  %��   	�  %��   	�k  %��   	�  %��   	Ӄ  %��   	�v  %��   	�a  %��   	�W  %��   	̶  %��   	�`  %��   	̨  %��   	��  %��   	��  %��   	��  %��   	�X  %��   	��  %��   	��  %��   	N�  &%T1  	��  &'�  �/  �8  	��  'My  	(h  'N�   	l�  'N�   	�  (.y  	�  (/y  	�  (0y  	�  (2y  	w�  (8�  	�  (9V  	�  (:�  	�_  (;�   	��  (>y  	�  (Jy  	"�  (R=  	t�  (S�   	�w  (T�   	؜  (Y�   	q�  ([y  	Ƚ  (^=  	�  (_�   	�y  (`�   	b�  (c�   	+�  (fy  	��  (iy  	֘ (l�   	�J  (x�   	��  (y�   	ks  (�   	�  (��   	J�  (��   	�i  (��   	��  (�y  	��  (�y  	��  (�y  	<� (�y  	��  (�y  	��  (�y  	5�  (�y  	<m  (��   	 K  (��   	�R  (��   	op  (��   	�m  (��   	D  (��   	X�  (��   	If  (��   	� (��   	��  (�y  	�U  (�y  	`  (�y  	J�  (�y  	��  (�y  	� (�p  -9  �O  =    	�  (��O  y  �O  =    	� (��O  U  �O  =   	 	,�  (��O  	R�  (��O  U  U  P  =    	�u  (��O  	��  (�R:  	�e  (��   �   CP  =   � 	(�  (�2P  	�  (�y  ��  (p  �v  (�   n�  (�   4�  (�   *b (�   ��  (M  	Y�  )%�%  	��  )&�%  	��  *.�  o	�P  x q	�    y q�    !�  r�P  t	Q  a v�P   b v�P   �u  w�P  y	EQ  x {8   y {8    �  |%Q  ~	qQ  a �EQ   b �EQ   ��  �QQ  �	�Q  slp �8   8{  �8   }  �}Q  qQ  �Q  =    +�e  �	�Q  	�^d     qQ  �Q  =    +�e  �	�Q  	�]d     qQ  	R  =    +[�  �	�Q  	@]d     +W�  �	�Q  	 ]d     ,k�  ��   	�e     ,)�  ��   	�e     -\�  ��   .�N  �	`�e     -W  ��   -�R  ��   /f_x ��   	 �e     /f_y ��   	��e     /f_w ��   	��e     /f_h ��   	��e     ,%]  ��   	�e     /fb ��  	�e     ,��  ��   	��e     ,�W  �EQ  	ؕe     ,�  �8  	Еe     ,`w  �8  	̕e     /m_x �8  	ȕe     /m_y �8  	ĕe     ,.�  �8  	��e     ,}  �8  	��e     /m_w �8  	��e     /m_h �8  	��e     ,��  �8  	��e     ,*x  �8  	��e     ,�  �8  	��e     ,�  �8  	��e     -y�  �8  ,A�  �8  	��e     -�c  �8  -,�  �8  ,�k  �8  	��e     ,�u  �8  	��e     ,�~  �8  	��e     ,^~  �8  	��e     ,a�  �8  	��e     ,�~  �8  	��e     ,�  �EQ  	��e     ,�k  �8  	�\d     0K\   8  	x�e     1plr  <  	p�e     M  vU  =   	 0"�  fU  	 �e     EQ  �U  =   	 0q^  �U  	��e     0q�  �   	��e     0��  �   	�\d     2�P  
	�\d     0�� y  	�\d     3�  :�%@     t       ��V  4�%@     _  BV  5U0 4&@     C[  ZV  5Uh 6&@     �Z  6&@     9X  4-&@     �W  �V  5Up5T@ 47&@     �V  �V  5Uu  6<&@     �V  7Z&@     �h   3'�  4�%@     %       ��V  8g  4�   U 3��  %@     �       ��W  9i !	�   |   z   9fx !�   �   �   9fy !�   �   �   9w !�   :  8  9h !�   `  ^  6A%@     �h  6k%@     �h  :�%@     �h  5Us   3��  �$@     d       �9X  ;��  �   �  �  ;wg  �   �  �  9i 
�       9t N1  |  z  :
%@     �X  5U	 ]d     5T35Q@@$  <��  ��X  =i �
�   =p � <  0��  �T1  	@KB     >g  �
�   >g  �
�    3~x  ��"@     �       �"Z  ;�  �"Z  �  �  ;��  ��   �  �  ;� �8      ;Mp ��  p  j  ;g  ��   �  �  ?x �8      @y �8  � 9i �
�   h  `  1l �qQ  ��44#@     �h  rY  5Uv  4C#@     �h  �Y  5Uv  4^#@     (Z  �Y  5U��5T��5Q|  4�#@     �h  �Y  5Uv  4�#@     �h  �Y  5Uv  4�#@     (Z  Z  5U��5T��5Q|  :�#@     \  5U��5T   qQ  3�c  �{"@     s       ��Z  ?x �j:  �  �  ?y �j:      ?a ��  o  k  A��  �8  �  �  6�"@     �h  4�"@     �h  �Z  5T~  4�"@     �h  �Z  5T~  6�"@     �h   3�h  c�!@     �       �C[  9i e	�   �  �  1l fqQ  	p�e     :q"@     \  5U	p�e       3�W  5� @     �       �\  ;g  5�   Q  K  9x 78  �  �  9y 78      A' 88  y  q  9end 88  �  �  1ml 9qQ  �P4%!@     \  �[  5Uw 5Tv  :�!@     \  5Uw 5Tv   3��  &� @             ��\  ?ml '"Z  =  9  ;g  (�   �  v  1fl *Q  	��e     4� @     �]  �\  5U�U5T	��e      B� @     �\  5U	��e     5T�T  3x�  ��@           ��]  ?fl ��]  	  
	  ;g  ��   b	  \	  9x ��   �	  �	  9y ��   �	  �	  9dx ��   �	  �	  1dy ��   P9sx ��   
  
  9sy ��   D
  B
  9ax ��   i
  g
  9ay ��   �
  �
  9d ��   �
  �
  0e  ��   	��e     B�@     �h  5T	2KB       Q  C`H  Py  �@     �      �_  ?ml Q"Z  �
  �
  ?fl R�]  t  j  !K   UU^  M �L 0�  )TOP  ATm  \�   �  �  Aʿ  ]�   �  �  A<�  ^�   7  5  9tmp `�P  l  Z  9dx a
�   r  V  9dy b
�   �  �  6L@     �h  6u@     �h  6�@     �h  6�@     �h   3�N  B�@            �;_  ;g  B�   �  �   3�  &O@     F       ��_  6m@     �_  6~@     B`  7�@     f   3x�  @     N       ��_  0�  �   	��e     0�  �/  	`KB     0�  �   	��e      3��  �.@     �       �B`  6f@     �h  6w@     �h  6�@     �h  :�@     �h  5Tv   3�G  ��@     R       ��`  6�@     �h  4 @     �h  �`  5U@<$ 7@     �b  7(@     lb  7.@     0g   C�d  Sy  �@     W      �Vb  ?ev TVb    �  9rc W	�   �  �  0�b  X�   	��e     0�< Y\b  	��e     9key Z	�   �  �  6�@     �b  4�@     �h  ca  5U@>$ 4#@     �h  |a  5U@>$ 4W@     �h  �a  5U@>$ 4�@     �h  �a  5U@>$ 6�@     zc  6@     g  6@     �b  6&@     �f  4�@     �h   b  5U	��e     5TD5Q	KB     5R	KB      6�@     �f  6	@     Ad  :;@     �h  5U	�\d         �   lb  =    3��  Gb@     #       ��b  4y@     �h  �b  5U@<$ 7�@     0g   3e�  =?@     #       ��b  4V@     �h  �b  5U@<$ 7b@     0g   3(P  *�@     ]       �zc  0Ī  ,�   	D\d     0�h  , �   	@\d     6�@     zc  6@     �c  69@     �e  7?@     �d   3�b  �@     &       ��c  0��    	P\d     6�@     td  :�@     i  5U	P\d       3�  G@     u       �Ad  6u@     Ad  6z@     0f  4�@     �h  +d  5T
3� :�@     �h  5U@<$  3;�  �&@     !       �td  9i �	�        36�  ��@     6       ��d  9i �	�   n  d  0��  �
rC  �g4@     i  �d  5U�g5T95Q	�JB     5Rs :@      i  5U�g  3�Y  ��@     E       ��e  9i �	�   �  �  0��  �
rC  �g4�@     i  me  5U�g5T95Q	�JB     5Rs  :�@     ,i  5U�g5T1  3�r  �f@     E      �f  AF� �	�   :  2  0��  �  	p\d     6�@     �h  6�@     �h  6z@     f  B�@     i  5U	p\d       D�t  ��@     �       �3��  c�@     +      ��f  9i e	�   �  �  9a f8      9b g8  >  <  6n@     �h  6�@     �h  :�@     �h  5T@A$  D��  W8@     J       �3�J  ?�@     �       �g  6@     �h  :0@     �h  5U@<$  D�  4X@     1       �3��  %�@     �       �jg  6�@     �h  6@     �h   3x�  ^@     ^       �h  ?ml "Z  e  a  ?is h  �  �  9dx 	�   �  �  9dy �       4�@     �h  �g  5Us 5Tv  :�@     �h  5Uv 5Ts   �Q  E9X  �#@     �       ��h  FGX  FRX  GtX  X  V  G�X    }  H�#@     X       �h  FGX  FRX  FtX  F�X  6=$@     �X   :�$@     �X  5U	�^d     5T75Q0  I��  ��  &EId  d  "	Iy�  y�  &9IF�  F�  bIH_  H_  #	IG�  G�  +/I�~  �~  3IY�  Y�  (	I[�  [�  fI�q  �q  $J	I��  ��  $C n3   �  S#  ]�  �*  	  2#  �)  �-   ,	  ^&  �  �1  @�   Q  �    �   	!   62  #	!     &	!   �5  )	!    �@  ,	!   (.  -	!   0*  2�   8;:  5�   < �   1  int �K 8"D   	�  K�   �   	�  L�   	�  M�   0t    e2    �0  }  ��    
;   Ji  D   �C  
D  ���� �C  NE  ڵ  R9  u  
;   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
;   /
  ��   [r  �4 #�  �   �X  5�  
;   :y  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K  
�   P�  =_  ��   R�  N�  ��  ��   �p  W�  
;   3�  ��   ({  ��  ğ   F]  8�  
;   Y0  ��   �c  |  ��  l  ��  �   
;   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {0  
;   ��  &�   �  º  GY  �f  ��   v�  ��  
;   �  GQ   ϼ  �  �_  X  &�  �b   
�	L  x �2   y �2  Mp �2  *� �2  ޽  �2   ~x �  	 	�  ��  	"+   E�  	#+  e% 	$2  u  	%
u  �8 	&
u  ��  	)
u  /b  	-
u  ��  	.	�   a  	2
u  �T  	3
u   Mx 	4X  �   �  �  	��  
Mi  	(h  
N�   	l�  
N�   	  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %'    �  -    	S�  '�  t�   �   �  �  �  -   �' �  	��  1�  	]  4�  �  �  �  -   � �  	Zy  8�  �  $  -   -   �   	��  ;$  Ʃ  Q;   5  A  W  -     F  	�  WW  �p  #�  S�  $�  �  �  B    T}  %�  �  �  B   B    '	�  acv )h  ��  *t  ��  +�   �y -�  �Y  6�  ��  :.  s�  <.   �H  =.  xz  >�   �  x @�  
;   �
  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �@  
;   �$$  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�
  (x	�$  �u z�
   � {	�   s |	�   � ~�  N�  $$  ��  �	�   ��  �	�     J]  �1$  �$  �$  -   � �^  ��$  �   �$    �  ��$  !;   �-(  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �$  \	�)  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /:(  �)  �)  -   � ��  1�)  
;   7�)  {�   U�  ~�   >	*  �� @*   s A
�   sx B�  sy C�   �$  Nz E�)  �]  ���+  `e �4   x ��  y ��  z ��   ��  ��+  (cN  ��+  0Mp �5  8�u ��
  <� ��   @�H  ��+  Hr�  ��+  P��  �,  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� �-(  �y� �,  �s ��   ��� �*  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  �+  ���  �   ���  	�   ��R  �-  �f�  �   �I}  L  ���  �+  �  *  "Gx  �+  �)  #d  HN�-  mo P'.   ��  Q.  cmd R�  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g-.  8�W  h=.  P��  ii  h�� lM.  l�N  m�  |E�  p�  ��W  r].  �~�  sM.  �*� tM.  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �'.  �$�R  ��    $��  ��   $�  ��   $h  �m.  $I�  �i  @ ,  �z  *  
;   1.  ��   ��  ��   �y  9�-  �-  �   =.  -    i  M.  -    �   ].  -    i  m.  -    *  }.  -    hy �,  (�	�.  in �i   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
M.  �a  �
�   $ ��  ��.  ��	�/  2�  �
�    I�  �i  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��/  ( �.  �/  -    ޴  ��.  	�  .i  	�  /i  	�  0i  	�  2i  	w�  8
  	�  9�  	�  :y  	�_  ;�   	��  >i  	�  Ji  	"�  R�  	t�  S�   	�w  T�   	؜  Y�   	q�  [i  	Ƚ  ^�  	�  _�   	�y  `�   	b�  c�   	+�  fi  	��  ii  	֘ l�   	�J  x�   	��  y�   	ks  �   	�  ��   	J�  ��   	�i  ��   	��  �i  	��  �i  	��  �i  	<� �i  	��  �i  	��  �i  	5�  �i  	<m  ��   	 K  ��   	�R  ��   	op  ��   	�m  ��   	D  ��   	X�  ��   	If  ��   	� ��   	��  �i  	�U  �i  	`  �i  	J�  �i  	��  �i  	� ��  }.  2  -    	�  �2  i  22  -    	� �"2  L  N2  -   	 	,�  �>2  	R�  �f2  L  L  |2  -    	�u  �l2  	��  ��/  	�e  ��   �   �2  -   � 	(�  ��2  	�  �i  ��  �  �v  �   n�  �   4�  �   *b �   ��  �  %�/  	�^d     %�/  	�e     %�/  	�^d     %0  	H-f     %0  		@-f      y    |  S#  h�  �*  �   &  ,   ,    2   1  Y�  %!   ��  &!   ,	  9   	@_d     E   #	 _d      �   �  S#  �  �*  [&@     d       �   G&  ,	  int ^&  9�  e2    �  �0  }  [   !�   �p   �  ��  S�  ��   �F  'p   *	�   *� ,�    "G  C	8   (G  C8   �]  C8   :G  C8    �U  D�   	�     
1   ? ��     	@�e     1�  8   	$�e     ��  8   	 �e     
�  +
�  �&@     2       ��  ��  -�  �  �   �   i�  #[&@     2       �ev #�  U  B%   �  S#  F�  �*  �#  (  �p  #-   3   :    S�  $F   L   W   W    T}  %e   k   {   W   W    	'	�   
acv )!   ��  *:   ��  +Y    �y -{       @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �  ��     ��  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u  (x	  �u z   � {	  s |	  � ~�   N�  �  ��  �	  ��  �	    int J]  ��  !  ?  ?  � ,	  �^  �.  ^  ^   d  1  �  �S    ��!  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � \	#  �Y  	   *O  	  ��  	  �  	  b�  	  ��  	  �  	  +�  	  Zp  	   o�   	  $m�  !	  (4�  "	  ,�  #	  0�  $	  4��  %	  8L� &	  <��  '	  @  (	  D��  )	  H\q *	  Lz�  +	  P�  ,	  T/�  -	  X ʤ  /�!  #  .#  ?  � ��  1#  �)  �?  ^&  �1  @�#  Q  ^   �   	;#  62  #	;#    &	;#  �5  )	;#   �@  ,	;#  (.  -	;#  0*  2  8;:  5  < �K 8"N#  �  K�#  �#  �  L�#  �  M�#  e2    �0  }    kt$  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
   ��$  &�   �  º  GY  �f  ��   v�  �t$  	%  ~�  �$   �S  
  ��   
    !
  �g  "
  �^  #
   ��  %�$  %  '%  ?   S�  '%  '%  %	�_d         R
  S#  E�  �*  �&@     �      v&  i)  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  9�  0t  4  e2    �0  }  ��  (  
K   J�  D   �C  
D  ���� �C  N\  ڵ  RP  
K   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
K   /  ��   [r  �4 #�  �   �X  5�  "	f  � $�    4h  %�  /  &  �_  '�     �  ((  f  	�  	�   	q  	�  �   	��  
%�   =� �  ��  .�  ^�  2o   }�  7u  �� ;K    	  r�  (   .� $9  O� )]   "  "  �    �    9  "   .  1   ]  "  K   R   1    ?  ��  ,�  c  �  oS  '�  dS  ()�  � +
�   � ,"  @�  -
�   >z .
�   �  /R   �H  3�    �   �  =    {  	�� 7�  	�� 8K   r  !  =      �  #!  	�PB     _�  <�  �   X  =    ��  =H  	`�e     ��  >�   	@�e     ��  A�   Y*@     5       ��  4h  A'�  U/  A;  Ti C	�   �  �   ��  2�   )*@     0       �.  4h  2'�  U/  2;  Ti 4	�        ��  �   *@     %       �t  �  (�  Ui 1   m  g   c�  �.  �)@     k       �.  � �#�   �  �  ��  �.    	  ��  �	�   `  X  ��  ��   �  �  i �	�   �)@     �    Ux �)@     V
  Uv �PB     "  4  r  ��  ��   �'@     �      ��	  � ��   �  �  4h  �+�	  &     ��  ��   �  r  1�  ��       ��  �	�   @  <  i �	�   |  v  �
  =(@     =(@     O       ��   �
  �  �   �
  �  �  !=(@     O       "
  *  (  "  R  N  ""  �  �  M(@     �  o  U} T/ v(@     �  U| Ts �PB     "   #.  �(@      P   �`	   Z  �  �   M  �  �   @  �  �  $P   "g  #    "t  \  Z  %�  �(@      �(@     }       � �  �  �   �  �  �  !�(@     }       "�  %    �(@     �  n  Uv T}  �(@     �  �  Uv  �(@     �  �  Uv  )@     �  �  Uv T	�XB      )@     �  �  U}  0)@     �  	  Uv T	(�B     Q} R0 B)@     �  0	  U	�NB     T}  J)@     �  H	  U}  V)@     �  U}      (@     �  �	  U	�NB     T1 &(@     V
  �	  Us  =(@       �	  U	�NB     Ts  �(@       �	  U	�NB      &�(@     �
   �  ��  ��   �'@            �V
  ��  � �   t  n  ��  ��   �  �  �'@     V
  Us   '��  t�   �
  (� t�   )�> v�   i w	�    *N�  7
'@     #       ��
  %G  
'@     
'@     "       h T  �  �    +P�  ��  .  (� �/�   (� �9�   i �1   )4h  ��  p ��    +��  ��   �  ,dir �+�   (� �4�   (4h  �I�	  )��  ��   i �1    +~�  ��   �  ,dir �*�   (�  �5�   )��  ��    -��  ��  �&@     K       �G  �> � �         ��  �,�   :   8   ��  �1   _   ]   `�  �1   �   �   �&@     �  T�T  .��  @a  /dir @�    0V
  -'@     �       ��   h
  �   �   1u
  1�
  2V
      t   h
  r!  j!  $    "u
  �!  �!  "�
  "  "  &L'@     �
  l'@     �  �  U} T|  x'@     �    U}  3�'@     �  �'@     �  F  T	(�B     Q| R0 �'@     �  ^  Uv  �'@     �  Uv    ?'@     �  Uv   4��  ��  A4��  ��  &4:�  :�  4$�  $�   	4��  ��  	4'�  '�  4��  ��  +4��  ��  d4m�  m�  @4��  ��  	%4��  ��  75      f   w  S#  ��  �*  �*@     q      P.  ,  �)  �=   ,	  int ^&  9�  0t  g   e2    �  �0  }  ��  [   u   J�   D   �C  
D  ���� �C  N�   ڵ  R�   u   K#  � � ^�  �� e  2 8� ��  �  _�  �   	�1  @�  
Q  �   
�   	1   
62  #	1   
  &	1   
�5  )	1    
�@  ,	1   (
.  -	1   0
*  2D   8
;:  5D   < �  1  �K 8"#  �  K�  �  �  L�  �  M�   	u  
��  "|    
E�  #|   
e% $�   
u  %
�   
�8 &
�   
��  )
�   
/b  -
�   
��  .	D   
a  2
�   
�T  3
�    Mx 4�  f 	�  �   �  =    g 
/�  	��  8
<  
{ 
@�   
x 
D�  
  
H�  
~  
N�  
1�  
R   
 �  
V  (
o  
Z(  0 R�  
0  	�   
4`  
"8 
6�   len 
71   
Q 
81   pos 
9u    i�  
1l  	��  
_�  
�> 
a.   
t 
bK    �   �   �  �  �  �   `    �  �   �  �  �   �  �  �    �  �  D    �    �     �  (  �     �  D
�	�  
w�  
�	D    
�  
�	D   
J�  
�	D   
�C  
�	D   
< 
�	D   
  
�	D   
� 
��  
��  
��  ,
5�  
�	D   @ I  
�4  d
�	�  
l�  
�	D    
n 
�	D   
֘ 
�	D   
K% 
�	D   
�  
�	D   
�  
�	D   
�  
�	D   map 
�	D   
  
�	D    
�  
�	D   $
J�  
�	D   (
\  
�	D   ,
b�  
�	D   0
:	 
�	D   4
 
�	D   8
�  
�	D   <
�R  
�	D   @
t 
�	�  D D   �  =    ��  
��  �   �  =    $
�	}  
�  
�	D    
� 
�	D   
 
�	D   
< 
�	D   
 
�	D   
�R  
�	D   
� 
�
}  ��  
�
}  � 
��  ���  
��    
�	D     �  �  =   =      
��  � �  �  �   �  D   D     	  
4 #
   
5# (&  
��  ,B  
|�  0
   
           D    u    <     <   �   ,  ! 1�  ��  M�   (h  ND   l�  ND   ��  ��  �\  ��   �  ��  �  ��  �D   ��  �D   2�  ��   ��  �D   Ɇ  ��  ��  �D   ��  �D   �h  �D   rK  �D   l�  �D   ]�  �D   ��  �D   �  D   q  K  �  t�   D   �C  %�   � &�   >�  '�  �  (�   � )�  �  +�  ��  ,�  2  -u   � .�  ��  /�  ��  0u   �C  2�   "�  `  � �  � �  � �  �-	A	  
��  /A	   
� 0�  � u  Q	  =    ��  1	  Q	  m	  =    � <]	  	��e     
 @D   	Пe     ��  DD   	̟e     `  H	P-f     T  		`�e     Z QD   @ UD   	ȟe     l  Z	\-f      ^Q  	T-f     \  b�   	X`d     7 fH
  	��e     H  � l�  	��e     5�  rD   	��e     ��  �
D   	X-f     � KD   	��e     D   �
  =    ��  L�
  	p�e     ��  MD   	h�e     � 7�/@            �   i 70H
  U � �--@     �      ��  !i �	D   �"  �"  "� �	D   �"  �"  "��  �	D   #  �"  / �D   	d�e     ")  �	D   e#  ]#  "��  �	D   �#  �#  "�} �	D   �$  �$  #@  �  !set �  %  %  $!  /@     p  0*  %/  S%  Q%  &p  '<  z%  v%  'I  �%  �%    (�  �/@     F       !l  )  *�/@     F       '  &  &    +�.@       �  ,U	/RB      -/@     �  ,Uv ,T~  .O/@     �  ._/@     U   $�  h-@     �   ��  &�   '�  �&  �&    /�  �-@     �-@     �       �A  *�-@     �       '�  �&  �&  '�  C'  ;'    $�  ~.@       o  &  '�  �'  �'    .=-@     "  .a-@     �  .h-@     �  .~.@     �  +�.@       �  ,U	RB      .�.@     "  +�.@     .  �  ,U1 .�.@     U   Q	  0��  �!  1set �-�  2i �u    0�  �U  1set �(�  2cmd �   2i �u    3� ��   �*@     ?       ��  "��  ��   �'  �'  !i �u   0(  .(   0 O�  2i Qu   4��  R	D    5  8D   �  4� :	D    6L 0�*@            �7Y �	�   -@             �j  8H �+j  Y(  S(  9��  ��    : -@     :  ,U	�*@     ,T1  �  t�  T�,@     :       ��  ;�  T)�  U;�� U0�  T �  !�  1�,@            ��  .�,@     �   U *,@     �       ��  8��     �(  �(  8��  /<  �(  �(  !i 	D   M)  I)  <�  :,@     �   	+K,@       r  ,U	�QB      =V,@     F  ,U	�QB        >� �?��  ��  J�  �	D   I �	D   @i �	D    Ab ��   �  ��  �	D   @cmd �u   Bl�  wD   �*@     .       �6  C[ y	D   �)  �)  .�*@     Q   D�  �*@     �       ��  '�  �)  �)  E�  Fm+@     T       �  E�  G�  �PH�+@     ,Uw   .+@     ]   I�  �+@     `       �  E�  E�  E�  &�   '�  *  *  '�  d*  Z*  '�  �*  �*  .�+@     �  .,@     �    J��  ��  7J  JB�  B�  !J  AK     J@ @ J� � � �s   �  S#  W �*  �/@     �      �7  �.  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  9�  0t  4  e2    �0  }  ��  (  
K   J�  D   �C  
D  ���� �C  N\  ڵ  RP  �  f �  �  �  =    	"|  *�  	��  +�  	I�  ,�  	�a  -�  
K   	4  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  	(�  
K   	/m  ��   [r  �4 #�  �   �X  	5@  
K   	:�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  	Ky  
�   	P  =_  ��   R�  N�  ��  ��   �p  	W�  
K   
3N  ��   ({  ��  ğ   F]  
8'  
K   
;�  �  � | 7	  �
 ` � � � 	 � 
FZ  
K   
Y�  ��   �c  |  ��  l  ��  �   
K   
k;  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  
{�  
K   
�z  &�   �  º  GY  �f  ��   v�  
�G  
K   
��  GQ   ϼ  �  �_  X  &�  �b   �   �  =    I  �  =    ;  �  =    
�	6  x �I   y �I  Mp �I  *� �I  ޽  �I   ~x ��   	�  ��  "B   E�  #B  e% $I  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4B  �  �   �  =    $�	�  �  �	�    � �	�    �	�   < �	�    �	�   �R  �	�   � �
�  ��  �
�  � ��  ���  ��    �	�     �   �  =   =      ��  �   �  �  	��  M�  	(h  N�   	l�  N�   	?  ~�  z   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�  ?  [  =    	S�  'K  t�   �   g  s  �  =   �' x  	��  1�  	]  4�  s  s  �  =   � �  	Zy  8�  �  �  =   =   � �  	��  ;�  Ʃ  QK   �      =       	�  W  �p  #�  S�  $@  F  Q  R    T}  %]  c  s  R   R    '	�  acv )(  ��  *4  ��  +Q   �y -s  �Y  6�  ��  :�  s�  <�   �H  =�  xz  >�   �  x @�  
K   Q  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  � 	  
K   ��%  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u]  (x	^&   �u zQ    � {	�    s |	�    � ~�   N�  �%   ��  �	�    ��  �	�     J]  ��%  ^&  |&  =   � !�^  �k&  �   �&  " !�  ��&  #K   ��)  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �&  \	G+   �Y  	�     *O  	�    ��  	�    �  	�    b�  	�    ��  	�    �  	�    +�  	�    Zp  	�     o�   	�   $ m�  !	�   ( 4�  "	�   , �  #	�   0 �  $	�   4 ��  %	�   8 L� &	�   < ��  '	�   @   (	�   D ��  )	�   H \q *	�   L z�  +	�   P �  ,	�   T /�  -	�   X ʤ  /�)  G+  d+  =   � !��  1T+  
K   7�+  {�   U�  ~�   >	�+  �� @�+   s A
�   sx Bg  sy Cg   ^&  Nz E�+  �]  ���-  `e ��   x �g  y �g  z �g   ��  ��-  (cN  ��-  0Mp ��  8�u �Q  <� ��   @�H  ��-  Hr�  ��-  P��  ��-  X��  �g  `m�  �g  d��  �g  h  �g  l3F  �g  p8F  �g  t=F  �g  x��  ��   |*� ��)  �y� ��-  �s ��   ��� ��+  ��  ��   ��  ��   �ʺ  ��   ��l  ��   �  �  �-  � ��  �   � ��  	�   � �R  �/  � f�  �   � I}  6  � ��  �-  � �+  Gx  ��-  >} �XE   �}  �I  �|  �I  
 �-  G+  $d  HN�/  mo P0   ��  Q0  cmd R�  �  Wg  (_  Yg   #_  [g  $bob ]g  (�  a�   ,�[  b�   0sb  d�   4d]  g0  8�W  h-0  P��  i�  h�� l=0  l�N  m;  |E�  p;  ��W  rM0  �~�  s=0  �*� t=0  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �0  ��R  ��    ��  ��   �  ��   h  �]0  I�  ��  @ �-  �z �+  
K   10  ��   ��  ��   �y  9�/  �/  �   -0  =    �  =0  =    �   M0  =    �  ]0  =    �+  m0  =    hy ��-  (�	�0  in ��   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
=0  �a  �
�   $ ��  �y0  ��	�1  2�  �
�    I�  ��  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��1  ( �0  �1  =    ޴  ��0  	�  .�  	�  /�  	�  0�  	�  2�  	w�  8m  	�  94  	�  :�  	�_  ;�   	��  >�  	�  J�  	"�  R  	t�  S�   	�w  T�   	؜  Y�   	q�  [�  	Ƚ  ^  	�  _�   	�y  `�   	b�  c�   	+�  f�  	��  i�  	֘ l�   	�J  x�   	��  y�   	ks  �   	�  ��   	J�  ��   	�i  ��   	��  ��  	��  ��  	��  ��  	<� ��  	��  ��  	��  ��  	5�  ��  	<m  ��   	 K  ��   	�R  ��   	op  ��   	�m  ��   	D  ��   	X�  ��   	If  ��   	� ��   	��  ��  	�U  ��  	`  ��  	J�  ��  	��  ��  	� �N  m0  4  =    	�  ��3  �  "4  =    	� �4  6  >4  =   	 	,�  �.4  	R�  �V4  6  6  l4  =    	�u  �\4  	��  ��1  	�e  ��   �   �4  =   � 	(�  ��4  	�  ��  !��  N  !�v  �   !n�  �   !4�  �   !*b �   !��  �  	Y�  %�&  	��  &�&  ) +5  J @�5  � "�    � '
�5  �� *	�   
 -�5  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 �   �5  =    5   H	6  � K�    C� N	�   "8 QR   t TR    . V�5  %6  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   5  u6  " 	R j6  6  �6  " 	� �6  
K   $E8  z  � �     & / 8 	; 
D M V _ h q z � q o z � � � � � � _ � o x �  � !�	 "  #1
 $� %< &( 'l
 (: )�	 *� +�
 ,� -V
 .# /� 0V 1� 2� 3� 4� 5a
 6� 7�
 8� 9� :D ;� <� =6 >f ?� @* Aa B C� D 
K   "�8  ��  WH  �~  �O  �m  ��   �  ��  ��  	 =� �8  ��  .�8  ^�  2X9   }�  7�  �� ;K    	�8  r�  9   .� $"9  O� )F9   &9  9  �    �8  �8  "9  9   9  &1   F9  9  K   R   1    (9  ��  ,�8  L9  oS  'j9  dS  ()�9  � +
�   � ,9  @�  -
�   >z .
�   �  /R   �H  3�9    ^9  	�� 7�9  	�� 8K   	 V�   	N�   %=0  	��   '�  
K   !!5:  �p   �  ��  S�  ��   �F  !':  !*	�:  *� !,5:   "G  !C	�   (G  !C�   �]  !C�   :G  !C�    �U  !DA:  
K   "�:  �  C	   	�  #�   	q  #�:  �   	��  $%�   	<]  %�   	��  %�   	h  %�   	��  %�   	�  %�   	�j  %�   	��  %�   	v  %�   	R  %�   	��  %�   	�o  % �   	�U  %"�   	�n  %#�   	�  %$�   	��  %%�   	�  %&�   	��  %'�   	u  %(�   	_b  %)�   	N  %*�   	�  %-�   	��  %.�   	0h  %/�   	�g  %0�   	��  %1�   	^�  %2�   	�a  %3�   	>�  %4�   	��  %5�   	O  %7�   	��  %8�   	Ϊ  %:�   	��  %;�  	ӄ  %=�   	r�  %>�   	~�  %?�   	��  %@�   	��  %A�   	��  %B�   	��  %C�   	��  %D�   	�T  %F�   		�  %G�   	^�  %H�   	��  %I�   	��  %J�   	�  %K�   	[n  %L�   	��  %M�   	-�  %O�   	��  %P�   	��  %Q�   	J�  %R�   	Ei  %T�   	��  %U�   	��  %V�   	A�  %W�   	��  %X�   	��  %Y�   	��  %Z�   	 t  %[�   	��  %\�   	!�  %]�   	oa  %^�   	/z  %_�   	��  %c�   	1P  %d�   	�  %e�   	Ʒ  %f�   	�T  %g�   	�o  %h�   	�b  %i�   	~�  %j�   	��  %k�   	�S  %m�   	��  %n�   	U  %o�   	Dl  %p�   	��  %q�   	��  %r�   	�p  %s�   	"�  %t�   	�  %u�   	�K  %v�   	��  %w�   	�  %y�   	tW  %z�   	'�  %{�   	��  %}�   	��  %~�   	�P  %�   	#L  %��   	gz  %��   	�  %��   	�k  %��   	�  %��   	Ӄ  %��   	�v  %��   	�a  %��   	�W  %��   	̶  %��   	�`  %��   	̨  %��   	��  %��   	��  %��   	��  %��   	�X  %��   	��  %��   	��  %��   	B &8�   	x	 &9�   	
 ':  	 ';�  w
 (6  	��  )��   	�\  )��  	�  )�_@  �  	��  )��   	��  )��   	2�  )��  	��  )��   	Ɇ  )��  	��  )��   	��  )��   	�h  )��   	rK  )��   	l�  )��   	]�  )��   	��  )��   	� *M�   	5 *N�   �   A  =   	 	~ +8A  H,#	�A  � ,'
�A   �^  ,(1    .�  ,)	�   (o�  ,-1   0i�  ,.	�   8��  ,/
�A  < �   �A  =    �   �A  =    �  ,0*A  	p�  -L�  	t�  -M�A  	K�  -N�A  	x�  -O�A  	��  -P�A  	��  -Q�A  	r�  -R�A  �A  B  =    	�  -SB  	�u  -T�A  		�  -U�A  	h�  -V�A  	��  ..�A  	�C  /%�  	� /&�  	>�  /'�  	�  /(�  	� /)�   	�  /+�  	��  /,�  	2  /-K   	� /.�  	��  //�  	��  /0K   	�C  /2�  C	�B  x Eg   y Fg   �{ H�B  (T	BC  `e V�   x Wg  y Xg  z Yg    	�  [
C  �a	(D  = cg   F�  dg  �~ eI  h�  fI  
t�  gI  �k hI  tag iI  �N  l
�   ��  o0  ��  r
=0   iK  uBC  0��  x
�   XS�  {0  `��  ~R   h��  ��   pu| ��D  x �}  X��D  v1 ��E   v2 ��E  dx �g  dy �g  �  �I  �k �I  tag �I  �W  ��  �o ��E  $��  ��E  4SX  �XE  8d�  �XE  @��  �
�   H��  �R   P �D  (D  �z �NC  �	XE  2�  �g   ]  �g  �h  �I  �N  �I  
�K  �I  >} �XE   �D  �}  � E  
K   ��E  ��   �  o�  ��   ��  �jE  �B  g  �E  =    �u  �(D  �z ��-  8�	;F  v1 ��E   v2 ��E  82  �g  Mp ��  [�  �;F   �  �AF   SX  �XE  (d�  �XE  0 ^E  �E  A{ ��E  4	�F  'x g   'y 	g  'dx 
g  'dy g   �o �F   )�  �  0 g  �F  =   =    (} SF  �  *�  (v  @2�G   @�  4�G   'x1 5�   'x2 6�    .]  8g   5]  9g   �� :g   ��  =�    �  @g    ��  Cg  $ �n  G�G  ( 9x  H�G  0 �^  I�G  8 GF  I  >�  K�F  (�h  PR�H   s�  U�H    �H  V�H  'x1 X�   'x2 Y�   'gx \g  'gy ]g  'gz `g   'gzt ag  $ �x  dg  ( � fg  , ~�  ig  0 t  kg  4 .� l�   8 �  p�H  @ 	�  r�   H �G  �F  �h  t�G  �	�H   �c  ��    �O  ��H   �x  �
�H   I  �H  =    �  �H  =    I�  ��H  �	(I   �  ��     �  �(I   �H  �  �I  )��	�I     �g    �  �	�    t�  �	�    ��  �	�    /�  �	�    �  �	�  'top �	�I  *��  �	�  U*��  �	�  V*� �	�I  W*�  �	�  � �  �I  =   ? ��  �;I  	.L  0&J  g  	׮  0)J  	�  0+J  	�  0,J  	�Q  0.�H  	��  00�   	��  01�   	(_  02�   	դ  04�   	�j  07�J  �   	��  08�J  	@�  0<�   	�O  0=�   	(g  0>�   	�^  0E�   	�u 0F�J  .I  	��  0H�   	��  0I�E  	��  0K�   	a� 0L�G  	w�  0N�   	P{ 0OXE  	��  0Q�   	��  0R5K  �E  	��  0T�   	�� 0USK  �F  	�}  0W�   	u| 0XAF  	M�  0Z�   	P�  0[;F  	��  0ag  	��  0bg  	�  0cg  	�p  0e�  	�T  0f�K  m0  	�a  0j�  �   �K  =   � 	ը  0l�K  �  L  =   @ 	�p  0m�K  	 �  0pg  	p|  0q�  	$Y  0v�   	�K  0y�   	g  0{ML  �I  	d�  0|ML  	��  1 g  		�  1!g  	�3 1#�   	_  1$�   	-�  1(�   	�f  1)�   	�G  1+g  	`�  1,g  	A�  1-g  	��  1/�   	��  11�   	P�  12�   �H  M  =   =   / 	��  1E�L  �H  !M  =   / 	Ԁ  1FM  �H  CM  =   =    	7� 1G-M  	�R  1I�   	��  1J�H  	��  1U�   	P�  1\6  	��  1]6  	L�  1^6  	ߵ  1_6  	�  1a6  	@�  2�G  	[�  2;F  	 �  2AF  	SX  2XE  	d�  2XE  	��  2�   	_�  2 �   	��  2"�  	��  2%�  	'�  2&�  	�]  2(�  �G  CN  =   � 	�P  2*3N  	ӯ  2+[N  �G  	|  2-mN  �H  	��  2.mN  	��  2/mN  �N  �N  �   �    	��  3�G  �  3 �N  	qY  3"�N  	�  3#�N  I  �N  =   ? 	��  3%�N  	��  3&�N  g  
O  =   � 	@Y  3(�N  g  'O  =   ? 	V�  3)O  �H  CO  =    	�h  43O  	�  4[O  �H  	�  4�H  	�f  4!�N  	r�  4"�N  	��  4%�G  	��  4&�G  	׆  4'g  	��  4(g  	�  4*g  	��  4+g  	�  5�H  	��  5�   	�_  5�   	�_  5�   	b  5g  	t  5g  	j�  5"�  	�  5:�   	��  5;�   	��  5<�   	�W  5>�H  	hn  5@g  	U~  5Ag  	�  5Bg  	 �  5Cg  	%�  5F�  	�u  5H�  	z  5I�  	� 6.�  +�4  Z	`6f     ,1�  ^�   	x-f     +�1  a
	`-f     -�1  b	d-f     -�1  c	,.f     -�1  d	$.f     	 j�  +2  l
	@2f     +"2  m	(.f     +.2  n	�-f     +F2  o
	�-f     +:2  p	D2f     ,� r
�  	0.f     ,a	 u�  	 .f     +�1  x	h-f     ,� {�  	��e     ,2�  }�4  	`2f     ,<
 ~�4  	@.f     ,� ��   	d`d     +�4  �	``d     	� ��  	*	 ��   .� ��   	l-f     .^ ��   	4.f     .f ��   	p-f     �   �R  =    /� \�R  �   �R  =    .�4 `�R  	�-f     �   �R  =    /� p�R  �S   �_  ��     � ��    �  ��   �R  /S  =   	 0� �S  	�\B     1�  �`:@     =	      �`  2p �	�   M+  %+  0� �
`  ��}0� �
�5  ��|35;@     �       T  4� 5
�   �,  �,  !��  6`  !E�  7`  5_;@     �n  6�;@     �n  7U	VB     7Ts   3�>@     \       �T  0� "`  ��|8i "�   9�>@     o  ]T  7U	�WB      9?@     o  uT  7Us  6)?@     o  7U	�WB       :�`  K<@       K<@            aU  ;a  2-  0-  <K<@            =a  9Z<@     �n   U  7U	WB     7Ts  6b<@     #o  7Us    >�`  n<@      @  k�U  ?@  @�`  ]-  U-  @�`  �-  �-  9}<@     /o  tU  7U	WB     7T1 9�<@     ;o  �U  7TsH�\B     " 9bC@     Go  �U  7U	�ZB      9C@     �n  �U  7U	WB      6�C@     o  7U	$WB        :�`  0>@      0>@     !       ��V  ;a  +.  !.  <0>@     !       @a  �.  �.  9D>@     �n  lV  7U	WB     7T��} 6Q>@     #o  7U��}   9y:@     Ro  �V  7U	.0@     7T0 9�:@     ^o  �V  7U	sUB      9�:@     Go  �V  7U	�UB      5�:@     jo  9�:@     vo  W  7U	�UB      9�:@     vo  0W  7U	�UB      9�:@     vo  OW  7U	�UB      9�:@     vo  nW  7U	�UB      5�:@     �o  9�:@     vo  �W  7U	�UB      9�:@     vo  �W  7U	�UB      9;@     Go  �W  7U	�UB      9#;@     �o  �W  7U0 9-;@     vo  X  7U	 VB      9�;@     Go  -X  7U	VB      5�;@     �o  9�;@     Go  YX  7U	4VB      9�;@     �o  �X  7U	nVB     7T	ZVB      5�;@     g  5�;@     �o  9<@     Ro  �X  7T0 9<@     �o  �X  7U? 90<@     o  �X  7U	zVB      9D<@     Go  Y  7U	�VB      9i<@     �o  #Y  7U0 5n<@     Fa  9�=@     o  OY  7U	>WB      9�=@     Go  nY  7U	GWB      5�=@     �o  9�=@     /o  �Y  7U	qWB     7T1 9�=@     /o  �Y  7U	{WB     7T1 9�=@     �o  �Y  7T	�WB      9>@     �o  Z  7U��}7Q
  90>@     �o  /Z  7U��}7T
 7Q	�WB      9�>@     �o  MZ  7U��|7Q9 9�>@     �n  sZ  7U	�WB     7T��} 9�>@     Ro  �Z  7T1 5�>@     p  5�>@     a  5�>@     p  5�>@     p  9<?@     o  �Z  7U	�WB      5E?@     *p  9O?@     Go  	[  7U	XB      9[?@     o  ([  7U	�XB      5k?@     6p  9u?@     o  T[  7U	�TB      9�?@     o  s[  7U	�TB      9�?@     Go  �[  7U	�XB      5�?@     *p  9�?@     Go  �[  7U	�YB      5�?@     Bp  5�?@     Np  5�?@     Zp  9�?@     fp  �[  7U1 5�?@     rp  5�?@     ~p  9�?@     /o  :\  7U	�YB     7T1 91@@     /o  ^\  7U	�YB     7T1 9|@@     /o  �\  7U	�YB     7T1 5�@@     �n  9�@@     vo  �\  7U	�YB      9�@@     /o  �\  7U	�YB     7T1 5�@@     �n  95A@     vo  �\  7U	>RB      9pA@     /o  "]  7U	�YB     7T1 5�A@     �n  9�A@     Go  N]  7U	�YB      5�A@     �p  9�A@     �n  z]  7U	�YB      5�A@     �p  9�A@     Go  �]  7U	ZB      5�A@     �p  9�A@     Go  �]  7U	3ZB      5�A@     �p  9�A@     Go  �]  7U	MZB      5 B@     �p  5B@     T`  9B@     Go  7^  7U	{ZB      5B@     �p  9B@     Go  c^  7U	�ZB      5#B@     �p  96B@     o  �^  7U	�ZB      9SB@     /o  �^  7U	�ZB     7T1 9fB@     Ro  �^  7T1 9pB@     Go  �^  7U	�ZB      9B@     /o  _  7U	�ZB     7T1 5�B@     �p  9�B@     /o  >_  7U	qWB     7T1 9�B@     �p  W_  7U��| 9�B@     /o  {_  7U	{WB     7T1 9�B@     �p  �_  7U��| 5�B@     �e  5�B@     q  9C@     �o  �_  7U��}7Q
  9C@     q  �_  7U��} 5JC@     q  5QC@     �d   �   `  =   � �   "`  =    �   8`  =   =    A )T`  /� +�   1i 7:@     )       ��`  2i 	�   �.  �.  B_:@     �n  7U	CUB       A� ��`  8p �	�   8i �	�    C3 ��`  8i �1   D/� ��     E�
 b�  a  F��  b �   /t d9   CE #Fa  /  %�  /� &�   1� ��7@     �      ��c  G   �a  8i �K   98@     &q  �a  7Us 7T	(TB     7Q8 9*8@     &q  �a  7UsX7T	.TB     7Q8 6F8@     o  7U	�TB       G@  �c  2p 	�   �.  �.  >�c  �8@       �  nc  ;�c  /  /  ?�  @�c  _/  M/  9�8@     2q  db  7Us 7T	CTB      9�8@     2q  �b  7Us 7T	ITB      9�8@     2q  �b  7Us 7T	MTB      99@     Go  �b  7U	VTB      9)9@     �n  �b  7U	oTB     7T	CTB      9:9@     �n  %c  7U	oTB     7T	ITB      9K9@     �n  Qc  7U	oTB     7T	MTB      B]9@     o  7U	tTB        6�8@     /o  7U	=TB     7T1  9\8@     o  �c  7U	3TB      6y8@     o  7U	8TB       A% �4d  F� �)�   8i �	�   �d   � ��     4h  ��    �c  0H �Dd  	�\B      d  Dd  =    4d  E ��   �d  FN � �   8i �1   /� ��   D/X �1   /�  ��     1� P�7@            ��d  HTe  �7@      �7@     
       T 1� �+6@     �      �Te  57@     >q  5u7@     �p  9�7@     2q  8e  7T	�SB      6�7@     o  7U	TB       I| �1� ��1@            ��e  9�1@     Jq  �e  7T8 B	2@     Vq  7U07T0  1� ��1@            ��e  HTe  �1@      �1@     
       � 1 �[5@     �       ��f  9�5@     Go  .f  7U	SB      5�5@     bq  5�5@     nq  5�5@     zq  5�5@     �q  9�5@     �q  �f  7U	�/@      5�5@     �q  5�5@     �q  5�5@     �q  5�5@     �q  5�5@     �q  5�5@     �q  5�5@     nq  56@     �q  56@     ji   JR �	�  1' O�0@     .      �Zi  2i Q	�   +0  #0  G�  �g  Kbuf wZi  �T9�1@     �q  �g  7U�T7T<7Q	�RB     7Rs 6�1@     �q  7U�T7Tvx  5�0@     
r  5�0@     r  5�0@     "r  5�0@     .r  5�0@     :r  5�0@     Fr  5�0@     Rr  5�0@     ^r  9�0@     jr  h  7U4 91@     �q  9h  7U	SRB      9(1@     �q  Xh  7U	eRB      971@     �q  wh  7U	pRB      9F1@     �q  �h  7U	}RB      9U1@     �q  �h  7U	�RB      9d1@     �q  �h  7U	�RB      9s1@     �q  �h  7U	�RB      9�1@     �q  i  7U	�RB      9�1@     �q  1i  7U	�RB      6�1@     �q  7U	�RB     7T	d`d       �   ji  =    L� �Nj  M� ��  	��e     MW ��  	��e     MS ��  	��e     MrK  ��  	��e     Mk	 �N  	\`d     M�	 ��   	��e     NJ�  ��   Ns ��   N� ��   Oy ��   N� ��  N ��  Nf ��   P2 �y0@     0       ��j  Qev ��j  �0  �0  5�0@     vr  9�0@     �r  �j  7Us  6�0@     �r  7Us   �:  R�f  �/@     /       �S8`  .0@     K       �yk  =F`  3X0@            ]k  @F`  �0  �0  9g0@     Jq  <k  7U	LRB     7T1 5o0@     �r  6v0@     �r  7U0  6T0@     vo  7U	>RB       Sji  	2@     R      �6n  =�i  =j  =j  =j  =)j  =5j  =Aj  ?�  @�i  1  �0  @j  ;1  71  @j  v1  r1  @j  �1  �1  @)j  �1  �1  @5j  2  2  @Aj  a2  [2  5-2@     �q  9b2@     �r  Ml  7U07T07Q
@7R� 5~2@     �r  5�2@     ^e  5�2@     �r  53@     �r  5(3@     �r  5/3@     �r  543@     �r  5T3@     s  5y3@     s  9�3@     Jq  �l  7U	�RB     7T8 5�3@     s  5�3@     *s  54@     6s  594@     Bs  9�4@     Jq  >m  7U	�RB     7T8 9�4@     Ns  Vm  7Tv  5�4@     Zs  5�4@     fs  T�4@     rs  9�4@     ~s  �m  7U07T07Q
@7R� 5�4@     �s  5�4@     �s  95@     �s  �m  7U1 9;5@     �s  n  7U17T07Q07R
@7X�7Y�\� 5C5@     �r  5H5@     Zs  5M5@     rs    RTe   6@            �Sa  a9@     �       ��n  @+a  �2  �2  @8a  �2  �2  G�  �n  =+a  =8a   9l9@     o  �n  7U	�TB      6x9@     o  7U	�TB       S�`  6:@            ��n  U�`    V� � 7(V��  ��  dV��  ��  (7Vj j <V� � :V��  ��  #%V'�  '�  8W    C V  (AVH H (MV� � 5V� � #!V# # )wV� � $V4 4  1V� � $"V� � $V��  ��  9,V� � LV�
 �
 :	V�	 �	 ;-	V  ;'	V[�  [�  fVZ Z E	V��  ��  9.VN N $#V	 	 (QV� � (IV� � )tVR R <$Vv v =?V� � �V�	 �	 �Vf f �V� � &0VC C 1�V� � >#V�
 �
  V	 	 �V� � +.VJ J -4V� � *4V( ( *(V� � *9V� � '#V� � *,V  *!V� � ?V:�  :�  ?Vn n =V��  ��  CVy�  y�   9VA A *6V� � >V� � )rV  )cV  )uV} } )aV� � )�V� �  VV�	 �	 �V!�  !�  AV� � )�V� � QVG�  G�  ;/V� � $V� � %�V� � )xV  =CV  �VC
 C
 %�Vg g %�V  %�V# # %�V  %�V
�  
�  !�
V e   e  &#	V�	 �	 *F	V� � @Vc� c� 7K#V� � "'V� � +6V�  �  .'V  -.VH H A(Vw w B%V�
 �
 )kV� � +4V� � 1�V� � )hV� � 5aVY Y 5dV�	 �	  iV� �  ?V�  �  &,V��  ��  7V  )lVG G "/V  <VB�  B�  <!V�
 �
 "7 S   �  S#  � �*  �C@     *      �K  �3  ,	  e2    �  �0  }  int ^&  F   J�   D   �C  
D  ���� �C  Ni   F   �   7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�   F   /  ��   [r  �4 #�  �   �X  5�   F   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K)  �  	4h  �    	/    	K% 	[   
map 	[    �  �  1    e  �  	�^B     w   	4h  x�    	�  y�   �  0  1   	 � z   	`^B     � �}  �D@            �}  4h  �)�   L3  H3   �  1  V �	�   �D@            ��  4h  �&�   U � �	�   eD@     3       �  4h  �*�   �3  �3  �  �A�  Ti �	[   �3  �3   � g[   8D@     -       ��  4h  g$�   �3  �3  /  g8  :4  44  K% i	[   �4  �4  WD@     �  Uu Tt Qy R1  � A	�   �C@     t       �	  4h  A)�   U/  A=  TK% B[   Qmap B,[   �4  �4  i D	[   =5  95   q 2	�   �C@     '       �4h  2'�   U/  2;  Ti 4	[   u5  s5    �=   T  S#   �*  �D@     �      �N  W4  �)  �=   ,	  int ^&  9�  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2D   8;:  5D   < �   1  �K 8"b   	�  K
  �   	�  L
  	�  M
  0t  4  e2    �0  }  ��  (  
[   J�  D   �C  
D  ���� �C  N\  ڵ  RP  �  
[   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
[   /!  ��   [r  �4 #�  �   �X  5�  
[   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K-  
D   P�  =_  ��   R�  N�  ��  ��   �p  W�  
[   3  ��   ({  ��  ğ   F]  8�  
[   ;Y  �  � | 7	  �
 ` � � � 	 � F  
[   Y�  ��   �c  |  ��  l  ��  �   
[   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {�  
[   �.  &�   �  º  GY  �f  ��   v�  ��  
[   �s  GQ   ϼ  �  �_  X  &�  �b   	� 	.Y  	�  
D   	q  
�  �   	B 8D   	x	 9D    	A  ��  "B   E�  #B  e% $I  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	D   a  2
�  �T  3
�   Mx 4�  �  	��  ��   	�\  ��  	�  �w  �  	��  �D   	��  �D   	2�  ��  	��  �D   	Ɇ  �M  	��  �D   	��  �D   	�h  �D   	rK  �D   	l�  �D   	]�  �D   	��  �D   	� MD   	5 ND   �   6  =    
�	}  x �I   y �I  Mp �I  *� �I  ޽  �I   ~x �6  f �  �  �  =    D�	$  w�  �	D    �  �	D   J�  �	D   �C  �	D   < �	D     �	D   � ��  ��  ��  ,5�  �	D   @ I  ��  d�	$  l�  �	D    n �	D   ֘ �	D   K% �	D   �  �	D   �  �	D   �  �	D   map �	D     �	D    �  �	D   $J�  �	D   (\  �	D   ,b�  �	D   0:	 �	D   4 �	D   8�  �	D   <�R  �	D   @t �	$  D D   4  =    ��  �0   	~  4 #�   5# (�  ��  ,�  |�  0�   �   ~  �  �  D    A  �  �  �  �   �  �  ! 1@  	��  M�  	(h  ND   	l�  ND   	K	  ~�  .   �S  
D   ��   
D     !
D   �g  "
D   �^  #
D    ��  %�  K	  g	  =    	S�  'W	  t�   D   s	  	  �	  =   �' �	  	��  1�	  	]  4�	  	  	  �	  =   � �	  	Zy  8�	  �  �	  =   =   � �	  	��  ;�	  Ʃ  Q[   
  
  #
  =     
  	�  W#
  �p  #�  S�  $L
  R
  ]
  K    T}  %i
  o
  
  K   K    '	�
  acv )4
  ��  *@
  ��  +]
   �y -
  �Y  6�
  ��  :�
  s�  <�
   �H  =�
  xz  >�
   �
  x @�
  
[   ]  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �  
[   ��'  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  ui  (x	j(  �u z]   � {	D   s |	D   � ~�
  N�  �'  ��  �	D   ��  �	D     J]  ��'  j(  �(  =   � �^  �w(  �   �(    �  ��(  ![   ��+  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �(  \	S-  �Y  	D    *O  	D   ��  	D   �  	D   b�  	D   ��  	D   �  	D   +�  	D   Zp  	D    o�   	D   $m�  !	D   (4�  "	D   ,�  #	D   0�  $	D   4��  %	D   8L� &	D   <��  '	D   @  (	D   D��  )	D   H\q *	D   Lz�  +	D   P�  ,	D   T/�  -	D   X ʤ  /,  S-  p-  =   � ��  1`-  
[   7�-  {�   U�  ~�   >	�-  �� @�-   s A
D   sx Bs	  sy Cs	   j(  Nz E�-  �]  ���/  `e �    x �s	  y �s	  z �s	   ��  ��/  (cN  ��/  0Mp �
  8�u �]  <� �D   @�H  ��/  Hr�  ��/  P��  ��/  X��  �s	  `m�  �s	  d��  �s	  h  �s	  l3F  �s	  p8F  �s	  t=F  �s	  x��  �D   |*� ��+  �y� ��/  �s �D   ��� ��-  ��  �D   ��  �D   �ʺ  �D   ��l  �D   � �  �/  ���  D   ���  	D   ��R  �1  �f�  D   �I}  }  ���  �/  � �-  "Gx  �/  S-  #d  HN�1  mo P�1   ��  Q�1  cmd RA  �  Ws	  (_  Ys	   #_  [s	  $bob ]s	  (�  aD   ,�[  bD   0sb  dD   4d]  g�1  8�W  h	2  P��  i�  h�� l2  l�N  m�  |E�  p�  ��W  r)2  �~�  s2  �*� t2  ��� wD   ���  xD   �X�  |D   ��e  D   ���  �D   �g  �D   ��u  �D   �|G ��   �Q  �D   ��  �D   �o�  ��1  �$�R  �D    $��  �D   $�  �D   $h  �92  $I�  ��  @ �/  �z �-  
[   1�1  ��   ��  ��   �y  9�1  �1  D   	2  =    �  2  =    D   )2  =    �  92  =    �-  I2  =    hy ��/  (�	�2  in ��   d  �
D   �x  �
D   D  �
D   5O  �
D   �� �
2  �a  �
D   $ ��  �U2  ��	^3  2�  �
D    I�  ��  r�  �
D   �H  �
D   *F  �
D   ��  �
D   	�  �
D   ѵ  �
D   ��  �
D    F� �
D   $�  �^3  ( �2  n3  =    ޴  ��2  	�  .�  	�  /�  	�  0�  	�  2�  	w�  8!  	�  9�  	�  :�  	�_  ;�   	��  >�  	�  J�  	"�  R�  	t�  SD   	�w  TD   	؜  YD   	q�  [�  	Ƚ  ^�  	�  _D   	�y  `D   	b�  cD   	+�  f�  	��  i�  	֘ lD   	�J  xD   	��  yD   	ks  D   	�  �D   	J�  �D   	�i  �D   	��  ��  	��  ��  	��  ��  	<� ��  	��  ��  	��  ��  	5�  ��  	<m  �D   	 K  �D   	�R  �D   	op  �D   	�m  �D   	D  �D   	X�  �D   	If  �D   	� �D   	��  ��  	�U  ��  	`  ��  	J�  ��  	��  ��  	� �  I2  �5  =    	�  ��5  �  �5  =    	� ��5  }  6  =   	 	,�  �
6  	R�  �26  }  }  H6  =    	�u  �86  	��  �n3  	�e  ��   �   }6  =   � 	(�  �l6  	�  ��  ��    �v  D   n�  D   4�  D   *b D   ��  �  =� �6  ��  .$7  ^�  2�7   }�  7M  �� ;[    	U7  r�  j7   .� ${7  O� )�7   %d7  d7  �    �6  U7  {7  d7   p7  %1   �7  d7  [   K   1    �7  ��  ,$7  �7  oS  '�7  dS  ()8  � +
&   � ,d7  @�  -
D   >z .
D   �  /K   �H  38    �7  	�� 78  	�� 8[   	"|  *�  	��  +�  	I�  ,�  	�a  -�  &�6  )	h6f     '2 a�  	�`d     (	 �WF@           �X:  '�  �4  ��)�;  xF@     �  �$9  *�;  �5  �5  +�F@     7=  9  ,U	�ZB      -�F@     7=  ,U	�_B       )�;  G@       �y9  *�;  �5  �5  .  /�;  6  �5  -�G@     C=  ,U	�_B        +xF@     N=  �9  ,U	�`d      +G@     Z=  �9  ,U��,T0 +�G@     f=  �9  ,U	2`B      +H@     f=  �9  ,U	q`B      +'H@     7=  :  ,U	�YB      +BH@     f=  2:  ,U	�`B      +UH@     r=  J:  ,Us 0_H@     C=   (f ��E@     �       ��;  'H �$  ��)�;  �E@      �  �\;  *�;  j6  f6  +�E@     7=  �:  ,U	�_B      +�E@     7=  �:  ,U	�_B      +�E@     7=  	;  ,U	�ZB      +F@     7=  (;  ,U	�_B      +F@     }=  @;  ,U�D -!F@     �=  ,U	�TB       +4F@     �=  u;  ,U�� -DF@     7=  ,U	�_B       1f ��;  2H �1�;   $  1F ��;  2�  �2�;   4  1� l�;  2�  l2�;  3i n[    4��  G�D@     �       ��<  5��  G�  �6  �6  5� G-�  �6  �6  	� I�  6i J[   I7  G7  )�<  �D@     p  R�<  7�<  .p  /=  o7  m7  +E@     �=  �<  ,U	 �e     ,T	�_B     ,QP 0VE@     �=    0uE@     �=  8�E@     �=   1W -!=  2�R  -&!=  ' /'=  	 �e     9� 0[    I2  �   7=  =   O :� � 
!;     :� � 4:t�  t�  J:��  ��  d;� �  :� �  :j j <:Y Y E	:  !'	:
 
 :	:� � 	':v v E 6Q   �  S#   �*  dH@     �
      JV  7  �  �)  �D   ,	  ^&  �1  @�   Q  �    �   	8   62  #	8     &	8   �5  )	8    �@  ,	8   (.  -	8   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
1   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �  	"|  *y  	��  +y  	I�  ,y  	�a  -y   	R  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�  
1   	!�  �p   �  ��  S�  ��   �F  	'^  	*	�  *� 	,�   "G  	C	�   (G  	C�   �]  	C�   :G  	C�    �U  	D�  
1   
"3  ��  WH  �~  �O  �m  ��   �  ��  ��  	 (	~  ��  B      B  Vd  !B  �  "B  �� #~   �   �  D    � %3  (	�  � *�   �� +�   � ,�  G /�  �   �  D    	N�  %�  	��  '�  �  �  
1   U  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (
  
1   /�  ��   [r  �4 #�  �   �X  5a  
1   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K�  
�   P<  =_  ��   R�  N�  ��  ��   �p  W	  =� T  ��  .�  ^�  2   }�  7�  �� ;1    	�  r�  �   .� $�  O� )   �  �  �    H  �  �  �   �  8     �  1   R   8    �  ��  ,�  
  oS  '(  dS  ()�  � +
�   � ,�  @�  -
�   >z .
�   �  /R   �H  3�    �   �  D      	�� 7�  	�� 81   t�   �   �  �  �  D   �' �  	��  1�  	]  4�  �  �    D   � �  	Zy  8  �  /  D   D   �   	��  ;/  Ʃ  Q1   @  L  b  D     Q  	�  Wb  �p  #  �  �   S�  $�  �  �  R    T}  %�  �  �  R   R    '	�  acv )s  ��  *�  ��  +�   �y -�  �Y  6�  ��  :F  s�  <F   �H  =F  xz  >     x @  
1   3  ��   ({  ��  ğ   F]  8X  
1   ;�  �  � | 7	  �
 ` � � � 	 � F�  
1   Y	  ��   �c  |  ��  l  ��  �   
1   kl	  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {	  
1   ��	  &�   �  º  GY  �f  ��   v�  �x	  
1   ��	  GQ   ϼ  �  �_  X  &�  �b   B   
  D    4  
  D    
�	W
  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x �
  
1   �  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �c
  
1   �G'  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�  (x	�'  �u z�   � {	�   s |	�   � ~�  N�  G'  ��  �	�   ��  �	�     J]  �T'  �'  �'  D   �  �^  ��'  �   �'  !  �  ��'  "1   �P+  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  (  \	�,  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /]+  �,  �,  D   �  ��  1�,  �]  ���.  `e �L   x ��  y ��  z ��   ��  ��.  (cN  ��.  0Mp �@  8�u ��  <� ��   @�H  ��.  Hr�  ��.  P��  ��.  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� �P+  �y� ��.  �s ��   ��� ��.  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  �.  ���  �   ���  	�   ��R  �0  �f�  �   �I}  W
  ���  �.  � �,  Gx  ��.  >} �+@   �}  �B  �|  �B  
 �.  �,  �'  #d  HN�0  mo P8   ��  Q
8  cmd RR  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g8  8�W  h,8  P��  iy  h�� l�  l�N  ml	  |E�  pl	  ��W  r<8  �~�  s�  �*� t�  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �8  �$�R  ��    $��  ��   $�  ��   $h  �L8  $I�  �y  @ �.  �z �,  ) �0  J @�1  � "�    � '
�1  �� *	�   
 -�1  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 �   �1  D    �0   H	�1  � K�    C� N	�   "8 QR   t TR    . V�1  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   �0  32  ! 	R (2  �1  J2  ! 	� ?2  
1   $4  z  � �     & / 8 	; 
D M V _ h q z � q o z � � � � � � _ � o x �  � !�	 "  #1
 $� %< &( 'l
 (: )�	 *� +�
 ,� -V
 .# /� 0V 1� 2� 3� 4� 5a
 6� 7�
 8� 9� :D ;� <� =6 >f ?� @* Aa B C� D 
1   r�6  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	 V�   	� .�  	Y�  %�'  	��  &�'  R  	��  My  	(h  N�   	l�  N�   	X7  ~�  �	   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  % 7  X7  t7  D    	S�  'd7  
1    7�7  {�   U�  ~�    >	�7  ��  @�.   s  A
�   sx  B�  sy  C�   Nz  E�7  
1   1
8  ��   ��  ��   �y  9�7  �0  �   ,8  D    y  <8  D    y  L8  D    �7  \8  D    hy ��.  (�	�8  in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�  �a  �
�   $ ��  �h8  ��	q9  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  �q9  ( �8  �9  D    ޴  ��8  	�  !.y  	�  !/y  	�  !0y  	�  !2y  	w�  !8�  	�  !9U  	�  !:�  	�_  !;�   	��  !>y  	�  !Jy  	"�  !R<  	t�  !S�   	�w  !T�   	؜  !Y�   	q�  ![y  	Ƚ  !^<  	�  !_�   	�y  !`�   	b�  !c�   	+�  !fy  	��  !iy  	֘ !l�   	�J  !x�   	��  !y�   	ks  !�   	�  !��   	J�  !��   	�i  !��   	��  !�y  	��  !�y  	��  !�y  	<� !�y  	��  !�y  	��  !�y  	5�  !�y  	<m  !��   	 K  !��   	�R  !��   	op  !��   	�m  !��   	D  !��   	X�  !��   	If  !��   	� !��   	��  !�y  	�U  !�y  	`  !�y  	J�  !�y  	��  !�y  	� !�  \8  �;  D    	�  !��;  y  <  D    	� !�<  W
  -<  D   	 	,�  !�<  	R�  !�E<  W
  W
  [<  D    	�u  !�K<  	��  !��9  	�e  !��   �   �<  D   � 	(�  !�<  	�  !�y   ��  !   �v  !�    n�  !�    4�  !�    *b !�    ��  !�6  	��  "��   	�\  "�y  	�  "�=  �  	��  "��   	��  "��   	2�  "�y  	��  "��   	Ɇ  "��  	��  "��   	��  "��   	�h  "��   	rK  "��   	l�  "��   	]�  "��   	��  "��   C	�=  x E�   y F�   �{ H�=  (T	>  `e VL   x W�  y X�  z Y�    	�  [�=  �a	�>  = c�   F�  d�  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  o8  ��  r
�   iK  u>  0��  x
�   XS�  {8  `��  ~R   h��  ��   pu| ��?  x �}  X��?  v1 �p@   v2 �p@  dx ��  dy ��  �  �B  �k �B  tag �B  �W  ��	  �o �v@  $��  �d@  4SX  �+@  8d�  �+@  @��  �
�   H��  �R   P �?  �>  �z �!>  �	+@  2�  ��   ]  ��  �h  �B  �N  �B  
�K  �B  >} �+@   �?  �}  ��?  
1   �d@  ��   �  o�  ��   ��  �=@  �=  �  �@  D    �u  ��>  �z ��.  8�	A  v1 �p@   v2 �p@  82  ��  Mp �@  [�  �A   �  �A   SX  �+@  (d�  �+@  0 1@  �@  A{ ��@  4	A  %x �   %y 	�  %dx 
�  %dy �  �o A  )�   
  0 �  �A  D   D    (} &A  �  *�  A  �A  �	�A  �c  �y   �O  ��A  �x  �
 B   B   B  D    �  B  D    I�  ��A  �	DB  �  ��    �  �DB   B  �  �B  &��	C    ��   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  %top �	C  '��  �	�  U'��  �	�  V'� �	C  W'�  �	�  � �  C  D   ? ��  �WB  	.L  #&+C  �  	׮  #)+C  	�  #++C  	�  #,+C  	�Q  #.�A  	��  #0�   	��  #1�   	(_  #2�   	դ  #4�   	�j  #7�C  �   	��  #8�C  	@�  #<�   	�O  #=�   	(g  #>�   	�^  #E�   	�u #F�C  JB  	��  #H�   	��  #Ip@  	��  #K�   	a� #L�A  	w�  #N�   	P{ #O+@  	��  #Q�   	��  #RQD  �@  	��  #T�   	�� #UoD  �A  	�}  #W�   	u| #XA  	M�  #Z�   	P�  #[A  	��  #a�  	��  #b�  	�  #c�  	�p  #e@  	�T  #f�D  \8  	�a  #j@  �   E  D   � 	ը  #l�D  @  !E  D   @ 	�p  #mE  	 �  #p�  	p|  #q@  	$Y  #v�   	�K  #y�   	g  #{iE  C  	d�  #|iE  
1   )�E  �  � 9  � -{E  (� 5�E  	�6f     (j 71   	�6f      <	F  4h  >U   K% ?	�   � ?�   U @�   � A�    � B�E  F  ;F  D    )� D+F  	�ad     (� a�   	�6f     (5 b�   	x6f     �   �F  D   	 	~ $8}F    �F  D   > 	D ��F  ,	�F  � .�    *� /P+   � 0�F  �F  �F  D    *� 2�F  	�`d     * H�   	�6f     *Z I�   	p6f     *q J
�.  	�6f     *� K
y  	�6f     *� L�   	�6f     *� M�   	�6f     *' N
y  	�6f     +w ��R@     x       �UH  ,UH  �R@     �  �:H  -�  .cH  �7  �7  / S@     qH  0<S@     �P   H  1T8 2IS@     �P  1U01T0   /�R@     AK  /�R@     �M   3{ �qH  4� ��    +R ^sQ@     _      �kJ  5� `�   �7  �7  6x a
�   #8  8  6p1 b  �8  �8  6p2 c  �8  �8  7� d
kJ  �V5� e
�   9  	9  7@ f�   	P�e     0�Q@     �P  @I  1U	�`B     1T5 0�Q@     �P  dI  1U	�`B     1T5 0�Q@     �P  �I  1U01T01Q
@1R� 0R@     {J  �I  1U| 0?R@     �P  �I  1U	�`B     1T8 0QR@     �P  �I  1Ul1TD 0�R@     �P  J  1U01T1 0�R@     �P  3J  1U�V1T:1Q	�`B     1Rs  0�R@     �P  PJ  1U�V1T8 8�R@     �P  1Ul1TD  �   {J  D   	 +� <Q@     V       �;K  9x =�   U:.� >  �9  �9  ;col ?�   �9  �9  5� A;K  :  	:  5m�  B�  6:  .:  5`5 C�  �:  �:  5� D�  *;  (;  5r� E
�   X;  R;   �  +d �P@     �       �YL  5� �C  �;  �;  5�  DB  �;  �;  5�O  !�   
<  <  5�x  "y  k<  g<  5.� #  �<  �<  0�P@     �P  �K  1U	�`B     1T8 0�P@     �P  	L  1U01T0 <�P@     YL  0 Q@     �P  -L  1T8 =Q@     	Q  KL  1U�1T� /Q@     �P   +� ��O@     �       �%M  :� ��   �<  �<  6ch ��   A=  7=  6c �
�   �=  �=  6cx �
�   B>  >>  6w �
�   z>  x>  5��  �
�   �>  �>  <.P@     Q  <\P@     Q  8�P@     �P  1Us 1T�  > �	y  DM  ?ev �#DM   �  @� f{M  Ast h
�   Asfx i
�   B+ � +� ToJ@     �       ��M  2�J@     !Q  1U?1T1  C� �dI@           ��N  Dsrc ��  �>  �>  E`5 ��  ?  ?  Dx �
�   �?  �?  Dy ��   �?  �?  Dw ��   �?  �?  Er� ��   E@  ?@  Dch ��   �@  �@  Dc �
�   �@  �@  Dcx �
�   @A  6A  Dcy �
�   �A  �A  0}I@     �P  �N  1T8 0�I@     �P  �N  1U01T01Q
@1R� <6J@     Q  8aJ@     �P  1U~ 1T|   C� ��N@     �       �MO  Fi �8   <�N@     {M  /�N@     JM  2NO@     -Q  1UN  GQ �	y  �O@            ��O  Hu �DM  �A  �A  2�O@     %M  1U�U  C ldH@            ��O  Fi n8   I�H@     �       �O  J{�  ��O   <�H@     !Q   F  KJM  �J@     �      �nP  LXM  LdM  -P  .XM  FB  >B  MdM  TNqM  �K@     0vK@     �P  YP  1U0 8�M@     �P  1U0   K%M  _O@     �       ��P  O7M  �B  �B  P%M  �  O7M  �B  �B  8�O@     �P  1U0   Q��  ��  CQy�  y�  9Q��  ��  EQ� � 6Q[�  [�  fQ� � BQ  :Q� � %QL L AQn n = �
   1   S#  Y �*  JS@     J      {b  �9  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"R   �  K  �   �  L  �  M  	K   "d  
��  
WH  
�~  
�O  
�m  
��  
 �  
��  
��  	 0t  p  e2    �0  }  ��  d  	K   J�  
D   
�C  
D  ���� �C  N�  ڵ  R�  �  ��  ��   �\  ��  �  ��  �  ��  ��   ��  ��   2�  ��  ��  ��   Ɇ  ��  ��  ��   ��  ��   �h  ��   rK  ��   l�  ��   ]�  ��   ��  ��   �   �  =    N�  	%�  ��  	'�  go #�  	x�e     2 %�  	p�e     � &�  	h�e     � '�  	`�e     y �(  	X�e     �   �
  �   �V@     �       �{   �   8C  4C  x �   uC  qC  y �   �C  �C  ��  �   �C  �C    �   CD  =D  G �   �D  �D  rc 	�   �D  �D  A 	{  	�B     ;W@       Uv T| Q}  IW@     �
  >  U0T0Qv R|  ]W@     ^  Uv T| Q}  �W@     Uv T| Q}   �  �  =    �  �   �  �   �   �    G ��   �V@     U       �q  x ��   E  E  y ��   ^E  XE  ��  ��   �E  �E    ��    F  �E  �V@     �
  ;  U
 �T1Q0 �V@     �
  �V@     �
  Us Tv Q| R�\�  � ��   |V@     %       �  x ��   ;F  7F  y ��   xF  tF  ��  ��   �F  �F    ��   �F  �F  �V@     �
    U
 �T1Q0 �V@     �
   { ��   �T@     )       ��  ��  ��   /G  +G    ��   lG  hG  G ��   �G  �G  U@     �
  U@     �
  U@     �
   M ��   �S@     4      �r  ��  ��   �G  �G     ��   TG ��   5H  1H  !i �
�   oH  kH  !j �
�   �H  �H  !dy �
�   ?I  ;I  !idx �
�   yI  uI  !s �r  �I  �I  !d �r  �J  �J  "� ��  �K  �K   �  � ��   �U@     �       �y  ��  ��   L  L    ��   jL  bL  G ��   �L  �L  !i �	�   M  M  !r ��   /M  -M  �U@     �	    T| Qs  �U@     �	  9  Tv 2Q�T V@     �
  ^  Uv 2$T1Qs  V@     �
  6V@     �
   � y�   �S@            ��   ��  z�   U   {�   T G |�   Q � K�   JS@     ^       �k	  ��  L�   `M  \M    M�   �M  �M   G N�   Q"� P�  �M  �M  !w Q�  \N  TN  !e R�  �N  �N  "� S
�   BO  >O   � A�   �T@            ��	  ��  B�   |O  xO    C�   �O  �O   G D�   Q #b +!U@     �       ��
  s ,
r  �O  �O  ��  -�   LP  DP    .�   �P  �P  !x 0
�   Q  �P  !y 1
�   ?Q  7Q  "`5 2r  �Q  �Q  GU@     �
  x
  Us T1Q0 $�U@     �
   %��  ��  	E%� � 6%  n%& & 	C%� � 7	%� � 
 x{   �"  S#  C  �*             �i  �;  �  int �)  �G   ,	  ^&  9�  �� �  �1  @�   Q  �    �   	;   62  #	;     &	;   �5  )	;    �@  ,	;   (.  -	;   0*  24   8;:  54   < �   1  �K 8"l   	�  K  �   	�  L  	�  M  0t  >  e2    �0  }  ��  2  
e   J�  D   �C  
D  ���� �C  Nf  ڵ  RZ  �  
e   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
e   /+  ��   [r  �4 #�  �   �X  5�  
e   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K7  
4   P�  =_  ��   R�  N�  ��  ��   �p  W�  
e   3  ��   ({  ��  ğ   F]  8�  
e   ;c  �  � | 7	  �
 ` � � � 	 � F  
e   Y�  ��   �c  |  ��  l  ��  �   
e   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {�  
e   �8  &�   �  º  GY  �f  ��   v�  �  
e   �}  GQ   ϼ  �  �_  X  &�  �b   �   �  G    S  �  G    E  �  G    
	�	�  x 	�S   y 	�S  Mp 	�S  *� 	�S  ޽  	�S   ~x 	��  
 	�  ��  
"L   E�  
#L  e% 
$S  u  
%
�  �8 
&
�  ��  
)
�  /b  
-
�  ��  
.	4   a  
2
�  �T  
3
�   Mx 
4   �  4   �  G    �   �  �  �  	��  M�  	(h  N4   	l�  N4   	C  ~�  8   �S  
4   ��   
4     !
4   �g  "
4   �^  #
4    ��  %�  C  _  G    	S�  'O  t�   4   k  w  �  G   �' |  	��  1�  	]  4�  w  w  �  G   � �  	Zy  8�  �  �  G   G   � �  	��  ;�  Ʃ  Qe   �      G     
  	�  W  �p  #�  S�  $D  J  U  N    T}  %a  g  w  N   N    '	�  acv ),  ��  *8  ��  +U   �y -w  �Y  6�  ��  :�  s�  <�   �H  =�  xz  >�   �  x @�  
e   U  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �  
e   ��$  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  ua  (x	b%  �u zU   � {	4   s |	4   � ~�  N�  �$  ��  �	4   ��  �	4     J]  ��$  b%  �%  G   � �^  �o%  �   �%    �  ��%  !e   ��(  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �%  \	K*  �Y  	4    *O  	4   ��  	4   �  	4   b�  	4   ��  	4   �  	4   +�  	4   Zp  	4    o�   	4   $m�  !	4   (4�  "	4   ,�  #	4   0�  $	4   4��  %	4   8L� &	4   <��  '	4   @  (	4   D��  )	4   H\q *	4   Lz�  +	4   P�  ,	4   T/�  -	4   X ʤ  /�(  K*  h*  G   � ��  1X*  
e   7�*  {�   U�  ~�   >	�*  �� @�*   s A
4   sx Bk  sy Ck   b%  Nz E�*  
e   p�+  �! 9& +! v( %# 0  B& @�! ��"  w#  	$  �-  S%  �)   0  @&  ��"    !0    m0    b-    �.    �$     /   @ %   � <"    U-    5'    	!  �]  ���-  `e ��   x �k  y �k  z �k   ��  ��-  (cN  ��-  0Mp ��  8�u �U  <� �4   @�H  ��-  Hr�  ��-  P��  ��-  X��  �k  `m�  �k  d��  �k  h  �k  l3F  �k  p8F  �k  t=F  �k  x��  �4   |*� ��(  �y� ��-  �s �4   ��� ��*  ��  �4   ��  �4   �ʺ  �4   ��l  �4   � �  �-  ���  4   ���  	4   ��R  �/  �f�  4   �I}  �  ���  �-  � �+  Gx  ��-  >} ��A   �}  �S  �|  �S  
 �-  K*  "d  HN�/  mo P�/   ��  Q�/  cmd R�  �  Wk  (_  Yk   #_  [k  $bob ]k  (�  a4   ,�[  b4   0sb  d4   4d]  g0  8�W  h0  P��  i�  h�� l!0  l�N  m�  |E�  p�  ��W  r10  �~�  s!0  �*� t!0  ��� w4   ���  x4   �X�  |4   ��e  4   ���  �4   �g  �4   ��u  �4   �|G ��   �Q  �4   ��  �4   �o�  ��/  �#�R  �4    #��  �4   #�  �4   #h  �A0  #I�  ��  @ �-  �z �+  
e   1�/  ��   ��  ��   �y  9�/  �/  4   0  G    �  !0  G    4   10  G    �  A0  G    �*  Q0  G    hy ��-  (�	�0  in ��   d  �
4   �x  �
4   D  �
4   5O  �
4   �� �
!0  �a  �
4   $ ��  �]0  ��	f1  2�  �
4    I�  ��  r�  �
4   �H  �
4   *F  �
4   ��  �
4   	�  �
4   ѵ  �
4   ��  �
4    F� �
4   $�  �f1  ( �0  v1  G    ޴  ��0  	�  .�  	�  /�  	�  0�  	�  2�  	w�  8+  	�  9�  	�  :�  	�_  ;�   	��  >�  	�  J�  	"�  R�  	t�  S4   	�w  T4   	؜  Y4   	q�  [�  	Ƚ  ^�  	�  _4   	�y  `4   	b�  c4   	+�  f�  	��  i�  	֘ l4   	�J  x4   	��  y4   	ks  4   	�  �4   	J�  �4   	�i  �4   	��  ��  	��  ��  	��  ��  	<� ��  	��  ��  	��  ��  	5�  ��  	<m  �4   	 K  �4   	�R  �4   	op  �4   	�m  �4   	D  �4   	X�  �4   	If  �4   	� �4   	��  ��  	�U  ��  	`  ��  	J�  ��  	��  ��  	� �  Q0  �3  G    	�  ��3  �  4  G    	� ��3  �  "4  G   	 	,�  �4  	R�  �:4  �  �  P4  G    	�u  �@4  	��  �v1  	�e  ��   �   �4  G   � 	(�  �t4  	�  ��  ��    �v  4   n�  4   4�  4   *b 4   ��  �  	"|  *�  	��  +�  	I�  ,�  	�a  -�  
e   "`5  ��  WH  �~  �O  �m  ��   �  ��  ��  	 
e   !�5  �p   �  ��  S�  ��   �F  '`5  *	�5  *� ,�5   "G  C	4   (G  C4   �]  C4   :G  C4    �U  D�5  
e   KA6  � � ^�  �� e  2 8� ��  �  _�  �   	�  4   	q  Y6  �   	<]  4   	��  4   	h  4   	��  4   	�  4   	�j  4   	��  4   	v  4   	R  4   	��  4   	�o   4   	�U  "4   	�n  #4   	�  $4   	��  %4   	�  &4   	��  '4   	u  (4   	_b  )4   	N  *4   	�  -4   	��  .4   	0h  /4   	�g  04   	��  14   	^�  24   	�a  34   	>�  44   	��  54   	O  74   	��  84   	Ϊ  :4   	��  ;�  	ӄ  =4   	r�  >4   	~�  ?4   	��  @4   	��  A4   	��  B4   	��  C4   	��  D4   	�T  F4   		�  G4   	^�  H4   	��  I4   	��  J4   	�  K4   	[n  L4   	��  M4   	-�  O4   	��  P4   	��  Q4   	J�  R4   	Ei  T4   	��  U4   	��  V4   	A�  W4   	��  X4   	��  Y4   	��  Z4   	 t  [4   	��  \4   	!�  ]4   	oa  ^4   	/z  _4   	��  c4   	1P  d4   	�  e4   	Ʒ  f4   	�T  g4   	�o  h4   	�b  i4   	~�  j4   	��  k4   	�S  m4   	��  n4   	U  o4   	Dl  p4   	��  q4   	��  r4   	�p  s4   	"�  t4   	�  u4   	�K  v4   	��  w4   	�  y4   	tW  z4   	'�  {4   	��  }4   	��  ~4   	�P  4   	#L  �4   	gz  �4   	�  �4   	�k  �4   	�  �4   	Ӄ  �4   	�v  �4   	�a  �4   	�W  �4   	̶  �4   	�`  �4   	̨  �4   	��  �4   	��  �4   	��  �4   	�X  �4   	��  �4   	��  �4   	B 84   	x	 94   �;  $	��  ��   	�\  ��  	�  �-   	��  �4   	��  �4   	2�  ��  	��  �4   	Ɇ  ��  	��  �4   	��  �4   	�h  �4   	rK  �4   	l�  �4   	]�  �4   	��  �4   	
 :  	 ;�  	� .c  �   �<  G   	 	~ 8r<  H #	�<  �  '
�<   �^   (;    .�   )	4   (o�   -;   0i�   .	4   8��   /
�<  < �   �<  G    �   =  G    �   0�<  	p�  !L�  	t�  !M=  	K�  !N=  	x�  !O=  	��  !P=  	��  !Q=  	r�  !R=  =  v=  G    	�  !Sf=  	�u  !T=  		�  !U=  	h�  !V=  	��  ".=  	N�  #%!0  	��  #'�  =� $�=  ��  $.>  ^�  $2�>   }�  $7�  �� $;e    $	<>  r� $ Q>   .� $$b>  O� $)�>   %K>  K>  �    �=  <>  b>  K>   W>  %;   �>  K>  e   N   ;    h>  ��  $,>  �>  oS  %'�>  dS  (%)?  � %+
}   � %,K>  @�  %-
4   >z %.
4   �  %/N   �H  %3?    �>  	�� %7?  	�� %8e   C	D?  x Ek   y Fk   �{ H$?  (T	�?  `e V�   x Wk  y Xk  z Yk    	�  [P?  �a	n@  = ck   F�  dk  �~ eS  h�  fS  
t�  gS  �k hS  tag iS  �N  l
4   ��  o�/  ��  r
!0   iK  u�?  0��  x
4   XS�  {�/  `��  ~N   h��  �4   pu| �.A  x �}  X�.A  v1 ��A   v2 ��A  dx �k  dy �k  �  �S  �k �S  tag �S  �W  ��  �o ��A  $��  ��A  4SX  ��A  8d�  ��A  @��  �
4   H��  �N   P 4A  n@  �z ��?  �	�A  2�  �k   ]  �k  �h  �S  �N  �S  
�K  �S  >} ��A   :A  �}  �FA  
e   ��A  ��   �  o�  ��   ��  ��A  D?  k  �A  G    �u  �n@  �z ��-  8�	�B  v1 ��A   v2 ��A  82  �k  Mp ��  [�  ��B   �  ��B   SX  ��A  (d�  ��A  0 �A  �A  A{ �B  4	�B  &x k   &y 	k  &dx 
k  &dy k  �o �B  )�  �  0 k  C  G   G    (} �B  �  *�  'v  @2�C  @�  4�C   &x1 54   &x2 64   .]  8k  5]  9k  �� :k  ��  =4   �  @k   ��  Ck  $�n  G�C  (9x  H�C  0�^  I�C  8 �B  S  >�  K"C  '�h  PR�D  s�  U�D   �H  V�D  &x1 X4   &x2 Y4   &gx \k  &gy ]k  &gz `k   &gzt ak  $�x  dk  (� fk  ,~�  ik  0t  kk  4.� l4   8�  p�D  @	�  r4   H �C  C  �h  t�C  �	E  �c  ��   �O  �E  �x  �
*E   S  *E  G    �  :E  G    I�  ��D  �	nE  �  �4    �  �nE   :E  �  �GE  (��	+F    �k   �  �	4   t�  �	4   ��  �	4   /�  �	4   �  �	�  &top �	+F  )��  �	�  U)��  �	�  V)� �	+F  W)�  �	�  � �  <F  G   ? ��  ��E  	.L  &&UF  k  	׮  &)UF  	�  &+UF  	�  &,UF  	�Q  &.�D  	��  &04   	��  &14   	(_  &24   	դ  &44   	�j  &7�F  4   	��  &8�F  	@�  &<4   	�O  &=4   	(g  &>4   	�^  &E4   	�u &FG  tE  	��  &H4   	��  &I�A  	��  &K4   	a� &L�C  	w�  &N4   	P{ &O�A  	��  &Q4   	��  &R{G  B  	��  &T4   	�� &U�G  C  	�}  &W4   	u| &X�B  	M�  &Z4   	P�  &[�B  	��  &ak  	��  &bk  	�  &ck  	�p  &e�  	�T  &fH  Q0  	�a  &j�  4   .H  G   � 	ը  &lH  �  KH  G   @ 	�p  &m:H  	 �  &pk  	p|  &q�  	$Y  &v4   	�K  &y4   	g  &{�H  <F  	d�  &|�H  	��  ' k  		�  '!k  	�3 '#4   	_  '$4   	-�  '(4   	�f  ')4   	�G  '+k  	`�  ',k  	A�  '-k  	��  '/4   	��  '14   	P�  '24   �D  KI  G   G   / 	��  'E5I  �D  gI  G   / 	Ԁ  'FWI  �D  �I  G   G    	7� 'GsI  	�R  'I4   	��  'J�D  	��  'U4   	P�  '\�;  	��  ']�;  	L�  '^�;  	ߵ  '_�;  	�  'a�;  	@�  (�C  	[�  (�B  	 �  (�B  	SX  (�A  	d�  (�A  	��  (4   	_�  ( 4   	��  ("�  	��  (%�  	'�  (&�  	�]  ((�  �C  �J  G   � 	�P  (*yJ  	ӯ  (+�J  �C  	|  (-�J  �D  	��  (.�J  	��  (/�J  �J  �J  4   4    	��  )�C  �  ) �J  	qY  )"�J  	�  )#�J  S  (K  G   ? 	��  )%K  	��  )&K  k  PK  G   � 	@Y  )(@K  k  mK  G   ? 	V�  ))\K  �D  �K  G    	�h  *yK  	�  *�K  �D  	�  *�D  	�f  *!K  	r�  *"K  	��  *%�C  	��  *&�C  	׆  *'k  	��  *(k  	�  **k  	��  *+k  	�  +�D  	��  +4   	�_  +4   	�_  +4   	b  +k  	t  +k  	j�  +"�  	�  +:4   	��  +;4   	��  +<4   	�W  +>�D  	hn  +@k  	U~  +Ak  	�  +Bk  	 �  +Ck  	%�  +F�  	�u  +H�  	z  +I�  	ʓ  ,C�  �  M  G    	��  ,b�L  4   #M  G    	��  ,cM  	0K  ,d4   	?�  ,e4   ,�	M  x ,�k   y ,�k  dx ,�k  dy ,�k   ��  ,�GM  ,��M  �p ,�
�/  ��  ,�
�B   ,�	�M  {q ,�k   ��  ,��  d ,�	�M   t�  ,��M  �M  �M  G   � 	r ,��M  	�T  ,�N  �M  	l�  ,�k  	�  ,�k  	?k  ,�k  	�d  ,�k  	2~ ,�M  	��  ,��  	��  ,�k  	k�  ,�k  	Z�  ,��B  �B  �N  G    	�v  ,��N  	�v  ,�4   	"�  ,��/  �  ,�  �U  ,�C  ��  ,�C  t�  ,4   �  ,	4   .Y  ,
k  7Y  ,k  �h  ,O  �/  *� ,!0  <i  ,!0  	G  -�  	��  -4   �   fO  G    
e   -��O  *top  �G  �  �]  -�fO   -�	�O  ��  -��B   ��  -��O  O{  -�
4   ��  -�
4   iK  -��O   �?  ��  -��O  �O   P  G    	��  -��O  !e   -3P  *up  �  �F  �S   FT  -
P  !e   -nP  ��   �x  H�  ��  �H   ��  -@P  H-	.Q  `e -�   >} -�A  L� -k   &low -k  $+� - k  (�Z -!
4   ,r� -"
4   0�f  -#3P  4�f  -$3P  8��  -%�  <&tag -&
4   @*� -'nP  D �w -){P  KQ  KQ  G    .Q  �  -2;Q  !e   -��Q  ��   �s  z�  ��  �T  ܭ   gY  -�^Q  H-�	6R  `e -��   *� -��Q  >} -��A   �W  -�k  (�}  -�k  ,L� -�k  0��  -��  4��  -�
4   8&tag -�
4   <��  -�
4   @  w -��Q  SR  SR  G    6R  j�  -CR  ) .rR  J @.S  � ."�    � .'
VO  �� .*	4   
 .-S  �9 .0	4    Ml  .3	4   $	
 .8	4   (C� .;	4   ,� .?	4   0� .BN   8 fR   .H	FS  � .K�    C� .N	4   "8 .QN   t .TN    . .VS  	: .�4   	3 .�4   	� .�4   	� .�4   	O .�4   	�
 .��   fR  �S    	R /�S  FS  �S    	� /�S  
e   /rkV  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	 0V4   	Y�  1%�%  	��  1&�%  	- 24   	_  2 4   	� 3M4   	5 3N4   +k	 ^  	49f     ,f<  `	89f     ,�3  a	09f     ,62  b	 Af     ,f2  c
	9f     ,B2  d	9f     ,N2  e	Af     ,Z2  i	 9f     -�2  k	�6f     +P! l�  	�;f     +�" m�  	9f     -�3  n	Af     +'- p�  	�7f     ,3  q	�;f     +�& r4   	p9f     ,3  t	�;f     ,~2  v	9f     -r2  w	�7f     ,4  x	�9f     -�3  y	�;f     + {�3  	�;f     ,>3  }	�6f     ,J3  ~	t9f     ,z3  	�;f     ,V3  �	X9f     ,b3  �	\9f     ,n3  �)	9f     +r% ��   	 9f     -�3  �	�;f     +	1 ��  	,9f     ,�3  �	x9f     -�3  �	�;f     + �
�  	(9f     +{0 ��  	P9f     +*1 ��  	@9f     ++ ��  	h9f     ,�3  �	H9f     ,�4  �	�ed     ,3  �	��e     ,&3  �	9f     ,\4  �	 Af     �  �Y  G   G    +��  ��Y  	�9f     k  Z  G    +��  ��Y  	�ed     +E�  ��Y  	�ed     k  CZ  G    +e% �3Z  	�ed     �F  iZ  G    .�" �YZ  	��B     .I- �4   	 �e     ��Z  ~�  ��   >- ��   �Z  �Z  �Z  G    �Z  .f' ��Z  	 �B     �  �Z  G   � .m1 ��Z  	 �e     .�  �4   	��e     .J/ �10  	��e     /~) ��  +�" �4   	�;f     +�" �4   	d9f     .1" �4   	��e     .2- ��  	��e     .A# �4   	��e     .% �4   	��e     .� ��  	��e     .& �4   	��e     .w/ �4   	��e     .� �4   	��e     .�& �4   	��e     �  I\  G    .�$ �9\  	@�e     /$ ��  .� �4   	 �e     �   �\  G    .m  ��\  	 �e     �/  �\  G    +�$ �
�\  	�6f     ,�4  �	`9f     ,�V  �	�ed     ,�V  �	�ed     4   ]  G   G   	 0r# ]  	 ed     4   @]  G    0q# !0]  	�dd     0E! -
�  	9f     f .�   � ��  �   �]  G   � 0W* �]  	 8f     0 �	�  	�;f     0I% �	4   	�9f     0�, �	4   	�;f     0o% 9�   	�;f     1
 �	�  �s@     X      �_  2�- �4   �Q  �Q  3�s@     K       �^  4fps �-   R  �Q  2)  �4   �R  �R  5�s@     %x  6�s@     1x  7U	��B       5�s@     =x  5et@     Ix  5lt@     Ux  5�t@     ax  5�t@     mx  6�t@     1x  7U	ÂB       8� �Is@     ;       �X_  9� ��   �R  �R  6Ws@     yx  7U	��B       8D' hNq@     �      �Ta  2  j�  3S  1S  4i k4   \S  VS  2K% k4   �S  �S  4map k!4   �S  �S  2�# l	4   �S  �S  3�q@     ^       �`  2|G ~�   T  T  :Ta  �q@      �q@     F       �	�`  ;fa  GT  ET  <�q@     F       6�q@     �x  7Uv 7T@7Q	��B     7Rs d7X	s d   5�q@     )b  6r@     �x  7U	��B     7Ts 7Rv   =mq@     �x  �`  7T1 5�q@     )b  =�r@     yx  a  7U	�_B      =s@     yx  "a  7U	��B      =s@     e  Fa  7Us 7Tv 7Q|  5*s@     %x   >' C�   �a  ?�  C)4   @�# E�a  	��e      �   �a  G    8( ;<q@            ��a  A� ;�   U 8A 
�o@     U      �)b  4i 4   nT  jT  =�o@     yx  b  7U	�_B      50p@     )b   1Q' �4   �o@     ?       �hb  6�o@     1x  7U	i�B       8� ��n@     �       �pc  9� ��   �T  �T  2�# �;   �T  �T  4i �	4   U  U  2�' �	4   -U  )U  =.o@     �x  �b  7Us 7T17Q0 =Oo@     �x   c  7Q	�WB     7Rv  =^o@     �x  Dc  7U	`�B     7T1 5uo@     �x  6�o@     �x  7Us 7T17Q0  8�/ �fu@     D      ��d  Bcmd �#�  rU  fU  2' ��  �U  �U  :�d  7v@      7v@     c       �Vd  <7v@     c       C�d  6V  4V  C�d  _V  YV  C�d  �V  �V  C�d  �V  �V  =Wv@     �x  Gd  7U~ 7T17Q0 5�v@     mx    5�u@     ^  D7v@     ^  E�v@     �d  7U�U  F2 ��d  G�& �	4   Gw0 ��  G9  ��  G� �	4    8� j�t@     �       �e  Bcmd j"�  *W  $W  D�t@     ^   8 ��k@     �      ��e  9  ��  ~W  vW  9K% �4   �W  �W  Bmap �4   �X  �X  2�) ��   Y  Y  4i �4   4Y  *Y  5�k@     �x  5^l@     �x  5�m@     �x  D�m@     s   8-  �un@     �       ��e  5�n@     e   8� ��k@            �@f  A  ��  UAK% �4   THmap �4   Q 8�, Jqj@     7      ��h  2� L�   �Y  �Y  2� M�   �Y  �Y  2�( N�   "Z  Z  5|j@     �x  5�j@     �x  =�j@     	y  �f  7Uv 7T	��B      =�j@     y  �f  7U	��B      =�j@     	y  !g  7Us 7T	��B      =�j@     1x  Lg  7U	��B     7Tv 7Qs  =�j@     !y  kg  7U	 �e      5�j@     -y  5�j@     9y  5�j@     Ey  5k@     Qy  5	k@     ]y  5k@     iy  =2k@     1x  �g  7U	ʀB      5>k@     uy  =Uk@     1x  h  7U	�B     7Tv 7Qs  =]k@     �y  (h  7U|  =hk@     �y  Fh  7Uv 7T|  =�k@     �y  xh  7U	 �e     7T	|�B     7Q  D�k@     �y   8�$ AOj@     "       ��h  9� B4   rZ  lZ  9�_  C	�   �Z  �Z  6ej@     �y  7U	 �e     7T�T7Q   I�/ i  G� 	4    8� 0j@            �ri  9� �   	[  [  6Cj@     �y  7U	 8f     7T�U7Q
   8�' ��i@     4       ��i  5j@     s   8�) ��i@     `       ��i  D�i@     �y   8q+ Bg@     }      �^j  4i D4   e[  U[  =@g@     �m  j  7Ux  5Wg@     �y  =�i@     �y  Bj  7U	 Af      E�i@     �y  7U	 Af       8�# 7�f@     A       ��j  6�f@     �y  7U	~�B       J�. 0�f@            �J�/ �f@            �I1 ��j  ?# �4   Ki �%4    8�% �ee@     �       ��k  9# �#4   \  \  4i �4   �\  �\  4j �4   �\  �\  2�' �4   ]  ]  =�e@     1x  �k  7U	Y�B     7T|  5�e@     �y  =�e@     �k  �k  7Us 7Tv  D�e@     �y   1�! \�  �c@     �      �Hm  9# ]4   V]  L]  9cp ^:4  �]  �]  4x `k  I^  G^  4y ak  n^  l^  4ss b{G  �^  �^  4mo c�/  �^  �^  4i d4   �^  �^  L`  �l  4xa �k  :_  ,_  4ya �k  �_  �_  4an �4   �`  t`  =e@     1x  �l  7U	7�B      64e@     z  7R'  = d@     z  m  7Ts 7Qv  5d@     z  =]d@     *z  3m  7Us 7Tv  6Xe@     6z  7T#  8�- 0�b@     �       ��m  9�R  04   �a  �a  4p 2H  �a  �a  4i 3
4   b  b  2�� 4
!0  �b  �b  2��  5
4   �b  �b  2g  6
4   c  c  2�u  7
4   uc  sc   8! ob@     V       �?n  9�R  4   �c  �c  4p H  �c  �c   8- �c@            ��n  9�R  4   @d  <d  E�c@     Hm  7U�U  8v V�v@     ;      ��p  4i X
4   �d  yd  4buf Y
4   Ee  9e  4cmd Z�  �e  �e  3�w@     B       Mo  @   ��p  	��e     � � q  6x@     �x  7U	��e     7TP7Q	�B       =�v@     �j  eo  7Us  5�v@     s  5w@     �e  5
w@     �h  5w@     @f  5w@     X_  5w@     �i  5&w@     �y  5-w@     ri  =9w@     Bz  �o  7U	ԂB      =�w@     �d  p  7U}  =�w@     pc  p  7U}  =�x@     1x  ;p  7U	��B      5y@     Nz  5y@     �x  =>y@     �y  �p  7U	 �e     7T	�B     7Q  5y@     Zz  D�y@     fz  5�y@     rz  5�y@     ~z  5�y@     �z  D�y@     �z  D�y@     �z  D�y@     �z   �    q  G   O �   q  G    1�	 �	�  �_@     �      ��r  Bev ��r  �e  �e  :�r  <a@       <a@     n       =	�q  ;�r  @f  >f  <<a@     n       C�r  if  cf  M�r  <a@     ]       C�r  �f  �f     :�r  �a@       �a@     l       C	5r  ;�r  �f  �f  <�a@     l       C�r  g  �f  Ms  �a@     [       Cs  Ug  Qg     5(`@     �z  =D`@     �z  Zr  7Us  =T`@     �z  rr  7Us  =d`@     �z  �r  7Us  6u`@     �z  7Us   �5  F�- ��r  ?� �*e   Ki �	4   NG�" �e     F�# �s  ?� �(e   Ki �	4   NG�" �4     8. [�]@     �      ��s  4i ]4   �g  �g  3^@     &       {s  2�) l�   �g  �g  5<^@     �x   =�]@     �z  �s  7U	�B      =�^@     {  �s  7Q0 5�^@     {   83# B�W@     Q      ��u  Bcmd B�  �g  �g  9
 B(4   Dh  @h  4i D
4   �h  }h  2R  E�  i  i  2��  F�  4i  2i  2L� G
4   Yi  Wi  2�. H
4   �i  |i  2�b  I
4   �i  �i  2<p J
4   %j  j  3�[@     *       �t  4key �4   �j  �j   3�]@             u  @�, FS  	��e     2]% GS  k  k   O�u  �Z@      �  �yu  ;�u  [k  Yk  P�  C�u  �k  ~k  Q�u  C�u  �k  �k  R�u  G[@          7;�u  �l  �l     5Z@     {   >�" 4   �u  ?��  4   G~�  �  G�& 	4   Ki 4    S�. ��  �u  T~�  �.�   U`* �4   �W@     	       �Av  Vcmd ��  UWi �;   �l  �l  Wsum �
4   Bm  8m   X�j  �e@     �       �w  ;�j  �m  �m  Q�j  Y�j  �  �v  ;�j  �n  }n  P�  C�j  o  �n  =\f@     �k  �v  7Us 7Tv  =uf@     �k  �v  7Us 7T}  =�f@     �y  �v  7U}  D�f@     �y    EDf@     �j  7U�U  X�h  �m@     �       �%x  Qi  L�  �w  Ci  So  Qo  5&n@     e  51n@     &{  56n@     2{  5;n@     >{  5@n@     J{  5En@     V{  =Sn@     1x  �w  7U	S�B      5_n@     uy  5mn@     b{  Dsn@     �y   =�m@     	y  
x  7U	 8f     7T	P�B      5�m@     o{  D	n@     uy   Z  4Z��  ��  57Z�q  �q  %J	Z/ / 55Z| | &Z�. �. 6	Z� � 7	Z� � !ZG�  G�  6/Z��  ��  dZ��  ��  %CZ� � 6Z��  ��  %Z� � 7(Z& & 0KZ�( �( 8$Zw! w! 90Z�/ �/ Z� � #Z�/ �/ [Z>1 >1 6ZE E (Z" " 1Z�( �( 3Z (  ( 5Z� � 7Z$ $ -ZpL pL �Z5L 5L YZ.' .' QZ�) �) RZ  6'	Z� � +aZ  :(Z�b  �b  "+Zm- m- ;Z�$ �$ <+Zj j %<Z� � 8![  YZ�( �( ,kZ�" �" ,�	Z11 11 ,qZ3, 3, '�Z� � 06Z3 3 #\Z$" $" 0JZ�) �) <.Z� � $Z�, �, =Ze$ e$ !+Z�  �  "#Z[$ [$ 3Z� � <$Z� � :"Z�  �  4Z,0 ,0 1	ZY�  Y�  !(	Z�d  �d  " 	ZQ Q :	Z) ) 9+Z8! 8! >Z[ [ ;	Z�. �. 5Zy' y' 2Z�) �) 4Z7. 7. 6Z�/ �/ 8Z�$ �$ ,	[�	 �	 �Z�& �& '	 >F   �'  S#  �3 �*  �y@     �      .�  �A  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �  
K   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {�  
K   �&  &�   �  º  GY  �f  ��   v�  ��  (	}  ��  B      B  Vd  !B  �  "B  �� #}   �   �  =    � %2  �   �  =    	N�  	%�  	��  	'�  �  �  t�  
 �   �  �p  #�  �  �   S�  $  	    R    T}  %   &  6  R   R    '	d  acv )�  ��  *�  ��  +   �y -6  �Y  6d  ��  :�  s�  <�   �H  =�  xz  >p   |  x @|  �  �  =   �' �  	��  1�  	]  4�  �  �    =   � �  	Zy  8  �  /  =   =   �   	��  ;/  Ʃ  QK   @  L  b  =     Q  	�  Wb  B  �  =    4  �  =    
�	�  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x ��  
K   7  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  
K   ��!  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  uC  (x	D"  �u z7   � {	�   s |	�   � ~d  N�  �!  ��  �	�   ��  �	�     J]  ��!  D"  b"  =   � �^  �Q"  �   z"   �  �o"   K   ��%  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �"  \	-'  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /�%  -'  J'  =   � ��  1:'  �]  ��-)  `e ��   x ��  y ��  z ��   ��  �-)  (cN  �-)  0Mp �@  8�u �7  <� ��   @�H  �-)  Hr�  �-)  P��  �h)  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� ��%  �y� �n)  �s ��   ��� �t)  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  -)  ���  �   ���  	�   ��R  T+  �f�  �   �I}  �  ���  -)  � W'  Gx  �h)  >} ��.   �}  �B  �|  �B  
 3)  -'  D"  !d  HNT+  mo Pl-   ��  Q�5  cmd R�5  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g
6  8�W  h6  P��  iy  h�� l�  l�N  m�  |E�  p�  ��W  r*6  �~�  s�  �*� t�  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �l-  �"�R  ��    "��  ��   "�  ��   "h  �:6  "I�  �y  @ z)  �z W'  	��  ��   	�\  �y  	�  ��+  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  ��  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	B,  x E�   y F�   �{ H",  (T	�,  `e V�   x W�  y X�  z Y�    	�  [N,  �a	l-  = c�   F�  d�  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  ol-  ��  r
�   iK  u�,  0��  x
�   XS�  {l-  `��  ~R   h��  ��   pu| �2.  x Z+  �}  X�2.  v1 ��.   v2 ��.  dx ��  dy ��  �  �B  �k �B  tag �B  �W  �s  �o ��.  $��  ��.  4SX  ��.  8d�  ��.  @��  �
�   H��  �R   P 8.  r-  �z ��,  �	�.  2�  ��   ]  ��  �h  �B  �N  �B  
�K  �B  >} ��.   >.  �}  �J.  
K   ��.  ��   �  o�  ��   ��  ��.  B,  �  �.  =    �u  �r-  �z �3)  8�	�/  v1 ��.   v2 ��.  82  ��  Mp �@  [�  ��/   �  ��/   SX  ��.  (d�  ��.  0 �.  �.  A{ �/  4	�/  #x �   #y 	�  #dx 
�  #dy �  �o �/  )�  �  0 �  0  =   =    (} �/  �  *�  $v  @2�0  @�  4�0   #x1 5�   #x2 6�   .]  8�  5]  9�  �� :�  ��  =�   �  @�   ��  C�  $�n  G�0  (9x  H�0  0�^  I�0  8 �/  B  >�  K&0  $�h  PR�1  s�  U�1   �H  V�1  #x1 X�   #x2 Y�   #gx \�  #gy ]�  #gz `�   #gzt a�  $�x  d�  (� f�  ,~�  i�  0t  k�  4.� l�   8�  p�1  @	�  r�   H �0  0  �h  t�0  �	2  �c  �y   �O  �2  �x  �
.2   B  .2  =    �  >2  =    I�  ��1  �	r2  �  ��    �  �r2   >2  �  �K2  %��	/3    ��   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  #top �	/3  &��  �	�  U&��  �	�  V&� �	/3  W&�  �	�  � �  @3  =   ? ��  ��2  p$	�3  x '
�    y (
�   f *�3  sc +
�   l ,
�3  len -
�   h�1 0
�   l �  �   �3  =   P �1 2M3  '�8	4  l :4   (h ;�   �(cl <�   �(on ?%4  �"R3 @y  � �3  %4  =    y  �2 B�3  �H	q4  l J�3   lm M�   pon P%4  xR3 Qy  � 2 S74  	�4  ~�  &   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %}4  �4  �4  =    	S�  '�4  >	95  �� @t)   s A
�   sx B�  sy C�   Nz E�4   	�5  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4E5  
K   1�5  ��   ��  ��   �y  9�5  �   6  =    y  *6  =    y  :6  =    95  J6  =    hy �z)  	.L  &b6  �  	׮  )b6  	�  +b6  	�  ,b6  	�Q  .�1  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�6  �   	��  8�6  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F"7  x2  	��  H�   	��  I�.  	��  K�   	a� L�0  	w�  N�   	P{ O�.  	��  Q�   	��  R�7  	/  	��  T�   	�� U�7  0  	�}  W�   	u| X�/  	M�  Z�   	P�  [�/  	��  a�  	��  b�  	�  c�  	�p  e@  	�T  f8  J6  	�a  j@  �   ;8  =   � 	ը  l*8  @  X8  =   @ 	�p  mG8  	 �  p�  	p|  q@  	$Y  v�   	�K  y�   	g  {�8  @3  	d�  |�8  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   �1  X9  =   =   / 	��  EB9  �1  t9  =   / 	Ԁ  Fd9  �1  �9  =   =    	7� G�9  	�R  I�   	��  J�1  	��  U�   )	P�  \�9  �9  	��  ]�9  	L�  ^�9  	ߵ  _�9  	�  a�9  	@�  �0  	[�  �/  	 �  �/  	SX  �.  	d�  �.  	��  �   	_�   �   	��  "y  	��  %y  	'�  &y  	�]  (y  �0  �:  =   � 	�P  *�:  	ӯ  +�:  �0  	|  -�:  �1  	��  .�:  	��  /�:  �:  �:  �   �    	��  �0  �   �:  	qY  ";  	�  #;  B  <;  =   ? 	��  %+;  	��  &+;  �  d;  =   � 	@Y  (T;  �  �;  =   ? 	V�  )p;  �1  �;  =    	�h  �;  	�  �;  �1  	�  �1  	�f  !+;  	r�  "+;  	��  %�0  	��  &�0  	׆  '�  	��  (�  	�  *�  	��  +�  	�  �1  	��  �   	�_  �   	�_  �   	b  �  	t  �  	j�  "�  	�  :�   	��  ;�   	��  <�   	�W  >�1  	hn  @�  	U~  A�  	�  B�  	 �  C�  	%�  F�  	�u  H�  	z  I�  	��  "y  *�2 T[~@     3       �S=  +it T#S=  |o  vo  ,�~@     wC  -Us   q4  *�1 IG~@            ��=  +it I"S=  �o  �o  .l L�=   p  p  /Z~@     D  -U�U-T1  �3  0�1 6y  ~@     ?       �Z>  +it 7S=  rp  lp  +ch 8-  �p  �p  1~@     F  '>  -U�T� 1(~@     �D  E>  -Us -Tt  ,6~@     W?  -Uu   *	3 *�}@     #       ��>  +it +S=  Sq  Oq  +str ,
�   �q  �q  ,�}@     �D  -Uu -Tt   *g3 #�}@            �?  2it ##S=  U3fE  �}@     �  &4sE  �q  �q    *�3 �}@            �W?  +it +S=  �q  �q  ,�}@     �D  -Uu   *�1 �}@            ��?  2it )S=  U/�}@     �D  -Uu   *=2 t}@     4       ��@  2it S=  U2x �   T2y 	�   Q5G 
�3  R5�1 �   X2on %4  Y3%E  �}@        4ZE  $r  "r  4PE  Ir  Gr  4FE  nr  lr  4<E  �r  �r  42E  �r  �r  6fE  �}@     `  ;4sE  �r  �r     7�2 �}@     U       ��@  8s �#�@  s   s  9i �	�   Xs  Rs  ,_}@     wC  -Uvps "  +4  7�2 ��|@     D       �gA  8s �"�@  �s  �s  9i �	�   �s  �s  9idx ��   It  Et  9l ��=  �t  �t  ,}@     D  -T0  7�2 ��|@     V       �B  8s ��@  �t  �t  :? �
�   u  	u  8msg �
�   Gu  Cu  1�|@     B  �A  -Uu  1�|@     �D  �A  -Uu -Tt  ,�|@     �D  -Uu -Tt   7�2 �+|@     Z       �|B  ;s �'�@  U9i �	�   �u  }u  <fE  M|@     M|@             �4sE  �u  �u    7�2 ��{@     l       �wC  8s ��@  v  v  ;x ��   T;y ��   Q;h ��   R=G ��3  X=�1 ��   Y;on �%4  � 9i �	�   [v  Uv  6%E  $|@      �  �4ZE  �v  �v  4PE  �v  �v  4FE  �v  �v  4<E  w  w  >2E  6fE  (|@     �  ;>sE     7>3 �{@     �       �D  8l �)�=  Fw  @w  9lh ��   �w  �w  9y ��   �w  �w  ?�2 ��   �w  �w  1�{@     )F  �C  -U|  @�{@     )F   7�1 ^dz@     �       ��D  8l _�=  x  x  :y1 `y  �x  �x  9i c�   	y  �x  9w d�   �y  {y  9x e�   �y  �y  9c f-  [z  Wz  @�z@     F  @�z@     5F  A{@     5F   B 2 P	y  Az@     #       ��D  ;t P2�=  U B%2 ?y  z@     *       �%E  ;t @�=  U;ch A
�   T C 3 0fE  Dt 1�=  Dx 2	�   Dy 3	�   Df 4�3  Dsc 5	�    Cs2 (~E  Dt ()�=   E33 $�y@            �FfE  �y@            ��E  GsE  U F%E  �y@            �F  G2E  UG<E  TGFE  QGPE  RGZE  X6fE  z@     @  ;4sE  �z  �z    H� � H�1 �1 6H� � 	? �M    ,  S#  �6 �*  �~@     �      l�  >D  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �  
K   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
K   /  ��   [r  �4 #�  �   �X  5�  
K   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K&  
�   P�  =_  ��   R�  N�  ��  ��   �p  W�  
K   3�  ��   ({  ��  ğ   F]  8�  
K   Y@  ��   �c  |  ��  l  ��  �   
K   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {@  
K   ��  &�   �  º  GY  �f  ��   v�  ��  
K   �  GQ   ϼ  �  �_  X  &�  �b   
K   	"Z  ��  WH  �~  �O  �m  ��   �  ��  ��  	 	"|  
*y  	��  
+y  	I�  
,y  	�a  
-y  �  	��  ��   	�\  �y  	�  ��  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  ��  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   
K   !x  �p   �  ��  S�  ��   �F  'K  *	�  *� ,x   "G  C	�   (G  C�   �]  C�   :G  C�    �U  D�  �   �  =   	 	~ 8�  t�   �   �  �p  #    !   S�  $-  3  >  R    T}  %J  P  `  R   R    '	�  acv )  ��  *!  ��  +>   �y -`  �Y  6�  ��  :�  s�  <�   �H  =�  xz  >�   �  x @�    �  =   �' �  	��  1�  	]  4      2  =   � !  	Zy  82  �  Y  =   =   � C  	��  ;Y  Ʃ  QK   j  v  �  =     {  	�  W�  �   �  =    B  �  =    
�	  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x ��  
K   a  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �  
K   ��$  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  um  (x	n%  �u za   � {	�   s |	�   � ~�  N�  �$  ��  �	�   ��  �	�     J]  �%  n%  �%  =   � �^  �{%  �   �%    �  ��%  !K   ��(  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �%  \	W*  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /
)  W*  t*  =   � ��  1d*  �]  ��W,  `e ��   x ��  y ��  z ��   ��  �W,  (cN  �W,  0Mp �j  8�u �a  <� ��   @�H  �W,  Hr�  �W,  P��  ��,  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� ��(  �y� ��,  �s ��   ��� ��,  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  W,  ���  �   ���  	�   ��R  ~.  �f�  �   �I}    ���  W,  � �*  Gx  ��,  >} �01   �}  �B  �|  �B  
 ],  W*  n%  "d  HN~.  mo PB0   ��  Q?  cmd R�=  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g$?  8�W  h4?  P��  iy  h�� lH0  l�N  m�  |E�  p�  ��W  rD?  �~�  sH0  �*� tH0  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �B0  �#�R  ��    #��  ��   #�  ��   #h  �T?  #I�  �y  @ �,  �z �*  (	�.  ��  B      B  Vd  !B  �  "B  �� #�.   �   �.  =    � %�.  C	/  x E�   y F�   �{ H�.  (T	\/  `e V�   x W�  y X�  z Y�    	�  [$/  �a	B0  = c�   F�  d�  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  oB0  ��  r
H0   iK  u\/  0��  x
�   XS�  {B0  `��  ~R   h��  ��   pu| �1  x �.  �   X0  =    �}  X�1  v1 �i1   v2 �i1  dx ��  dy ��  �  �B  �k �B  tag �B  �W  ��  �o �o1  $��  �]1  4SX  �01  8d�  �01  @��  �
�   H��  �R   P 1  X0  �z �h/  $1  
K   �]1  ��   �  o�  ��   ��  �61  /  �  1  =    p$	�1  x '
�    y (
�   f *�1  sc +
�   l ,
�1  len -
�   h�1 0
�   l �1  �.  �   �1  =   P �1 21  $�8	M2  l :M2   %h ;�   �%cl <�   �%on ?]2  �#R3 @y  � �1  ]2  =    y  �2 B2  �H	�2  l J�1   lm M�   pon P]2  xR3 Qy  � 2 So2  	<]  �   	��  �   	h  �   	��  �   	�  �   	�j  �   	��  �   	v  �   	R  �   	��  �   	�o   �   	�U  "�   	�n  #�   	�  $�   	��  %�   	�  &�   	��  '�   	u  (�   	_b  )�   	N  *�   	�  -�   	��  .�   	0h  /�   	�g  0�   	��  1�   	^�  2�   	�a  3�   	>�  4�   	��  5�   	O  7�   	��  8�   	Ϊ  :�   	��  ;�.  	ӄ  =�   	r�  >�   	~�  ?�   	��  @�   	��  A�   	��  B�   	��  C�   	��  D�   	�T  F�   		�  G�   	^�  H�   	��  I�   	��  J�   	�  K�   	[n  L�   	��  M�   	-�  O�   	��  P�   	��  Q�   	J�  R�   	Ei  T�   	��  U�   	��  V�   	A�  W�   	��  X�   	��  Y�   	��  Z�   	 t  [�   	��  \�   	!�  ]�   	oa  ^�   	/z  _�   	��  c�   	1P  d�   	�  e�   	Ʒ  f�   	�T  g�   	�o  h�   	�b  i�   	~�  j�   	��  k�   	�S  m�   	��  n�   	U  o�   	Dl  p�   	��  q�   	��  r�   	�p  s�   	"�  t�   	�  u�   	�K  v�   	��  w�   	�  y�   	tW  z�   	'�  {�   	��  }�   	��  ~�   	�P  �   	#L  ��   	gz  ��   	�  ��   	�k  ��   	�  ��   	Ӄ  ��   	�v  ��   	�a  ��   	�W  ��   	̶  ��   	�`  ��   	̨  ��   	��  ��   	��  ��   	��  ��   	�X  ��   	��  ��   	��  ��   =� �7  ��  .8  ^�  2�8   }�  7�  �� ;K    	C8  r�  X8   .� $i8  O� )�8   &R8  R8  �    �7  C8  i8  R8   ^8  &1   �8  R8  K   R   1    o8  ��  ,8  �8  oS  '�8  dS  ()9  � +
�   � ,R8  @�  -
�   >z .
�   �  /R   �H  39    �8  	�� 79  	�� 8K   ) 79  J @�9  � "�    � '
�9  �� *	�   
 -�9  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 �   �9  =    +9   H	:  � K�    C� N	�   "8 QR   t TR    . V�9  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   +9  z:    	R o:  :  �:    	� �:  
K   r@=  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	 V�    	�=  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4L=  �=  	��  My  	(h  N�   	l�  N�    	f>  ~�   �   �S   
�   ��    
�      !
�   �g   "
�   �^   #
�    ��   %>  f>  �>  =    	S�   'r>  
K   !7�>  {�   U�  ~�   !>	�>  �� !@�,   s !A
�   sx !B�  sy !C�   Nz !E�>  
K   1?  ��   ��  ��   �y  9�>  �   4?  =    y  D?  =    y  T?  =    �>  d?  =    hy ��,  (�	�?  in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
H0  �a  �
�   $ ��  �p?  ��	y@  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  �y@  ( �?  �@  =    ޴  ��?  	�  ".y  	�  "/y  	�  "0y  	�  "2y  	w�  "8  	�  "9�  	�  ":�  	�_  ";�   	��  ">y  	�  "Jy  	"�  "R�  	t�  "S�   	�w  "T�   	؜  "Y�   	q�  "[y  	Ƚ  "^�  	�  "_�   	�y  "`�   	b�  "c�   	+�  "fy  	��  "iy  	֘ "l�   	�J  "x�   	��  "y�   	ks  "�   	�  "��   	J�  "��   	�i  "��   	��  "�y  	��  "�y  	��  "�y  	<� "�y  	��  "�y  	��  "�y  	5�  "�y  	<m  "��   	 K  "��   	�R  "��   	op  "��   	�m  "��   	D  "��   	X�  "��   	If  "��   	� "��   	��  "�y  	�U  "�y  	`  "�y  	J�  "�y  	��  "�y  	� "��  d?  �B  =    	�  "��B  y  C  =    	� "�	C    5C  =   	 	,�  "�%C  	R�  "�MC      cC  =    	�u  "�SC  	��  "��@  	�e  "��   �   �C  =   � 	(�  "��C  	�  "�y  ��  "�  �v  "�   n�  "�   4�  "�   *b "�   ��  "�=  	Y�  #%�%  	��  #&�%  '�  @	�jd     �   8D  =    (� N(D  	`jd     (�4 V�   	Df     )plr WzD  	p�e     d?  �1  �D  =   > (D X�D  	 Bf     *�4 Y�1  	 �e     (�5 Zy  	Bf     *e5 [�2  	`�e     *s5 \y  	D�e     �   E  =    *[5 ]�D  	@�e     �2  4E  =    *�5 ^$E  	 �e     *�4 `y  	�e     (�5 ay  	 Bf     *A5 by  	�e     *�6 dc2  	@�e     *15 e�   	$�e     	*	 g�   *#5 iy  	 �e     �   �E  =   , (�5 p�E  	�hd     �   F  =   _ (�4 � F  	�ed     �   6F  =    +�5 �&F  	��e     +�  ��   	��e     +�W ��   	|�e     ,,0  	y  ��@     �      �`H  -ev  `H  �z  �z  +�6 �1  	 �e     .56 �   �{  z{  .l5 y  �{  �{  +5 y  	x�e     /c -  �|  �|  /i �   ,}  }  .�5 	�   �}  �}  +5 �   	t�e     0{�@     �L  {G  1U	`�e      2��@     �H  0 �@     �L  �G  1U	`�e      2��@     �H  0��@     �H  �G  1Uu  0�@     �L  �G  1U	 �e     1QQ 0
�@     M  H  1U	`�e     1Tv � 0�@     �H  1H  1Uu  3F�@     �L  1U	 �e     1T	t�e     1QQ  �  ,�. ��   ˂@     %       ��H  /c �
�   ~  ~   4�4 ���@     6       ��H  5c ��   U 4[$ �ۀ@     �      ��I  /i �	�   ?~  ;~  /rc ��   y~  w~  /c �
�   �~  �~  0G�@     M  GI  1U	@�e     1T0 0�@     M  hI  1U~ 1T| � 07�@     M  �I  1U	@�e     1Qv 4�e     " 0o�@     M  �I  1U0 3w�@     �L  1U~   4� ���@             �<J  0ƀ@     'M  J  1U	@�e      0Ѐ@     3M   J  1U	`�e      6ۀ@     ?M  1U	 �e       4� ��@     -       ��J  0��@     KM  zJ  1U	@�e      0��@     WM  �J  1U	`�e      6��@     cM  1U	 �e     1T0  4�4 4�~@     �      �+L  7i 7
�   /s 8�   �~  �~  8+L  �~@     �~@     
       ;0]@     oM  ZK  1U	@�e     1T01Q01R11X	 Bf     1Y! 0�@     {M  �K  1U	 �e     1T01R	 Bf     1X! 0'�@     �M  �K  1U	 �e      0]�@     �M  �K  1U	`�e     1T01R	 Bf     1X!1Y	Bf      3{�@     �M  1Us�~1T01Q01R01X01Y	D�e       9�3 /4� �~@     F       ��L  /i !
�     �~  /j "
�   S  M  +�< #
�9  �g0�~@     �M  �L  1U�g1T91Q	ĄB     1Rs! 3�~@     �M  1U�g1T1  :+L  �~@            �;g3 g3 �;  $'	;�1 �1 �;�2 �2 �;� � 6;�2 �2 �;�2 �2 �;>3 >3 p;�2 �2 �;�1 �1 �;�1 �1 m;�2 �2 y; 3  3 d;%2 %2 g	;=2 =2 �;[�  [�  f;��  ��  C =*   ~/  S#  �6 �*  ��  �G  �)  �-   ,	  ^&  �  �1  @�   Q  �    �   	!   62  #	!     &	!   �5  )	!    �@  ,	!   (.  -	!   0*  2�   8;:  5�   < �   1  int �K 8"D   	�  K�   �   	�  L�   	�  M�   9�  0t  $  e2    �0  }  ��    ڵ  R@  
L  ) i  J @�  � "�    � '
�  �� *	�   
 -	  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BB   8 �   	  -    ]   H	M  � K�    C� N	�   "8 QB   t TB    . V  d  B    Y  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   ]  �   	R �  M  �   	� �  ;   r�  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m t�   �   
�  �p  	#�  �  �   S�  	$d  T}  	%�  �  �  B   B    	'		  acv 	)�  ��  	*�  ��  	+�   �y 	-�  ;   
f	  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  
�  ;   
��"  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  
ur	  (
x	s#  �u 
zf	   � 
{	�   s 
|	�   � 
~	  N�  
�"  ��  
�	�   ��  
�	�     J]  
�#  s#  �#  -   � �^  
��#  �   �#   �  
��#  ;   
�'  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � \
	O(  �Y  
	�    *O  
	�   ��  
	�   �  
	�   b�  
	�   ��  
	�   �  
	�   +�  
	�   Zp  
	�    o�  
 	�   $m�  
!	�   (4�  
"	�   ,�  
#	�   0�  
$	�   4��  
%	�   8L� 
&	�   <��  
'	�   @  
(	�   D��  
)	�   H\q 
*	�   Lz�  
+	�   P�  
,	�   T/�  
-	�   X ʤ  
/'  O(  l(  -   � ��  
1\(  �  �(  -   �' 
y(  	��  1�(  	]  4�(  �  �  �(  -   � 
�(  	Zy  8�(  X  �(  -   -   � 
�(  	��  ;�(  Ʃ  Q;   
�(  )  )  -     
)  	�  W)  ;   p	*  �! 9& +! v( %# 0  B& @�! ��"  w#  	$  �-  S%  �)   0  @&  ��"    !0    m0    b-    �.    �$     /   @ %   � <"    U-    5'    	!   �#   	@3e      �#  		 �d     !l(  J	�jd      O   1  S#  �7 �*          #       l�  aI  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"R   �  K  �   �  L  �  M  e2    �0  }  �6 �   	;  $	        
Y7 ��   v  �7 ��    
8 ��   �7 ��   z7 ��                  ��  Ml  ��   U l7 ��   �7 ��   �7 k�   �  �6 k�    7 \               �7 &�                    ��                 ��  U  v   y2  S#  ?8 �*  p�@            ?�  �J  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"R   �  K  �   �  L  �  M  0t  +  e2    �0  }  ��    	K   Jw  
D   
�C  
D  ���� �C  NS  ڵ  RG  �  ��  ��   �\  �w  �  ��  �  ��  ��   ��  ��   2�  �w  ��  ��   Ɇ  ��  ��  ��   ��  ��   �h  ��   rK  ��   l�  ��   ]�  ��   ��  ��   � $p�@            �8 $�  U  n   C3  S#  9 �*  q�@     �       �  �K  �)  �=   ,	  int ^&  9�  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2D   8;:  5D   < �   1  �K 8"`   �  K  �   �  L  �  M  e2    �0  }  ��  %�   	J8 0D   	��e     	�8 4D   	�7e     	�8 9D   	��e     	�8 :D   	��e     	�8 ?D   	�7e     	�8 @D   	|�e     	i8 DD   	�7e     	�8 ED   	x�e     
D     =   	 	~8 I�  	�7e      St�@     �       �  i U	D   �  �  �  �  � b  �@�@     Y  �  Uw T Q	�B     Rs  �@     e  Uw Tv|  ��@     e  �  U	v�B     T	��e      ��@     e    U	��B     T	�7e      ��@     e  ?  U	��B     T	��e      ��@     e  k  U	��B     T	�7e      ̅@     e  �  U	��B     T	�7e      ۅ@     e  �  U	ǓB     T	��e      �@     e  �  U	ٓB     T	|�e      ��@     e  U	�B     T	x�e       
�   (  =    %9 Av sV8 M1  r�@            �G�  G�  /� �  .+   �4  S#  �9 �*          �      ǫ  �M  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"R   �  K  �   �  L  �  M  9�  0t  2  e2    �0  }  ��  &  	K   J~  
D   
�C  
D  ���� �C  NZ  ڵ  RN   (	�  ��  ,	�      -	�   &: 4�  �9 9  �= Y~   �  �   �  �  ~    �   �   �   �    �  ]< Z�  ��  ��   �\  �~  �  �L  �  ��  ��   ��  ��   2�  �~  ��  ��   Ɇ  ��  ��  ��   ��  ��   �h  ��   rK  ��   l�  ��   ]�  ��   ��  ��   �  �   q  �  �   	K   	"F  
��  
WH  
�~  
�O  
�m  
��  
 �  
��  
��  	 �< %�  	        z: )�  	        D: -�   	        �  �  =    &= 4�  	        >< 8�  	        : `  	        O: �  	        k: �  	        �: �  	        ]:   	        K; �  	        �; e  	        �; �  	        �; �  	        < �  	        �: ?  	        ; �  	        <; �  	        r; d  	        �; �  	        g; �~  �  x1 ��   y1 �'�   x2 �/�   y2 �7�   �: ��  e9 ��  y �	�    /: n�  `5 n.�  src n:�  x p	�   c q	�   M9 r�  S9 r�  Y9 r�  _9 r#�   1; J~  \  x1 J�   y1 J'�   x2 J/�   y2 J7�   �: L�  e9 L�  y M	�    �< ��  `5 �.�  src �:�  x 	�   c 	�   M9 �  S9 �  Y9 �   ; �~  *  x1 ��   y1 �'�   x2 �/�   y2 �7�   �: ��  e9 ��  y �	�    �9 ��  `5 �.�  src �:�  M9 ��  S9 ��  x �	�   c ��    �: �~  �  x1 ��   y1 �'�   x2 �/�   y2 �7�   �: ��  e9 ��  y �	�    �9 N7  `5 N.�  src N:�  M9 P�  x Q	�   c Q�    �: %~  �  x1 %�   y1 %'�   x2 %/�   y2 %7�   �: '�  e9 '�  y (	�    �9 �  `5 .�  src :�  x 	�    k< �~  ;	  x1 � �   y1 �(�   x2 �0�   y2 �8�   �: ��  e9 ��  y �	�    �; �        +       ��	  `5 �&�  �  �  src �2�  _�  Y�  x �	�     Q< ~  �	  x1  �   y1 (�   x2 0�   y2 8�   �: �  e9 �  y 	�    ;         9       ��
  `5 -�  ��  ��  �; 9�  /�  '�  �; E�  ��  ��  C< &�  R x 		�   �  �   val 
	�   e�  c�   [; �        #       ��
  `5 �&�  ��  ��  src �2�  �  
�   x �	�   ��  �   2< �~  T  x1 � �   y1 �(�   x2 �0�   y2 �8�   �: ��  e9 ��  y �	�    �< z        2       ��  `5 z-�  ׃  у  �; z9�  (�  "�  �; zE�  ��  }�  C< {&�  R x }	�   ܄  ؄   val ~	�   �  �   : l        !       �G  `5 l&�  C�  =�  src l2�  ��  ��   x n	�   �  �   �; ~  �  x1  �   y1 (�   x2 0�   y2 8�   �: �  e9 �  y 	�    �:         /       �E  `5 -�  ,�  $�  �; 9�  ��  ��  �; E�  �  �  C< 	&�  R x 	�   ��  ��   val 	�   ߇  ݇   �: �               ��  `5 �&�  �  �  src �2�  ��  ��   x �	�   ��  ��   �; �~  
  x1 � �   y1 �(�   x2 �0�   y2 �8�   �: ��  e9 ��  y �	�    �: �        )       ��  `5 �-�  S�  K�  �; �9�  ȉ  ��  �; �E�  =�  5�  C< �&�  R x �	�   ��  ��   !m9 �        �       �z  @� ��  �  ��  "        �*  "        �*  #        �*  �  $U	         #        �    $Us $TD #        �  3  $Us $T( "        �*  #        �*  _  $U	         %        �  $Us $T2  ;9 ��  @� �%�   �: i�  @� i'�   &< L�          L      �S  @� L)�  T�  N�  pct L6�   ��  ��  '��  N�  ��  ��   x O	�   ]�  [�   y O�   ��  ��   r P	�   �  ݌   g P�   �  �   b P�   Y�  U�  '69 Q�  ��  ��  '�9 R�  э  ͍  (S          �  _#3  )�  �  	�  )}  G�  E�  )r  n�  l�  )e  ��  ��  *�  +�  ��  ��  +�  ��  �  +�  5�  /�  +�  ��  ��  +�  ď      %        �*  $U@<$$T1$Q0  �; '�   �  @� '#�  r '0�   g '7�   b '>�   col )�  < *	�   �< +	�   �< ,	�   i -	�    ,�9 �~          �      �n  -x1 ��   �  �  -y1 �&�   (�  $�  .x2 �.�   Q-y2 �6�   e�  a�  /�: ��  ��  ��  /e9 ��  ǐ  ��  /�= ��  �  �  /�= �'�  i�  _�  /�; �2�  ��  ��  /�= �=�  i�  a�  0x �	�   В  ̒  0y ��   �  �  /�9 �	�   A�  =�  *�   sp  �  ��  ��   sp2  �  f�  X�   sp3  �  6�  (�   sp4   �  �  ��   sp5  &�  ֖  Ȗ   bp  ,�  ��  ��    ,�< �~          �       ��  .x1 ��   U-y1 �&�   �  �  .x2 �.�   Q.y2 �6�   R/�: ��  (�  &�  /e9 ��  M�  K�  /�= ��  r�  p�  /�= �'�  ��  ��  /�; �2�  ��  ��  0x �	�   �  ߘ  0y ��   k�  i�  /�9 �	�   ��  ��  *�  0sp ��  ��  �  0sp2 ��  ֚  Ț  0sp3 ��  ��  ��  0sp4 � �  ��  ��  0bp �&�  j�  b�    ,w< �~          �       �  -x1 ��   �  ��  -y1 �&�   !�  �  .x2 �.�   Q.y2 �6�   R/�: ��  \�  Z�  /e9 ��  ��  �  /�= ��  ��  ��  /�= �'�  ˞  ɞ  0x �	�   �  �  0y ��   <�  :�  /�9 �	�   e�  _�  *@  0sp ��  ş  ��  0sp2 ��  ]�  S�  0sp3 ��  ��  �  0bp � �  ��  ��    ,�9 i~          �       �  .x1 i�   U-y1 i&�   ء  ԡ  .x2 i.�   Q.y2 i6�   R/�: k�  �  �  /e9 k�  <�  6�  /�= k�  ��  ��  0x l	�   ڢ  ΢  0y l�   x�  r�  /�9 m	�   ǣ  ã  *   0sp v�  �  ��  0sp2 v�  ��  ��  0bp v�  I�  A�    ,�9 K~          _       ��  -x1 K�   å  ��  -y1 K&�    �  ��  -x2 K.�   =�  9�  -y2 K6�   z�  v�  /�: M�  ��  ��  /e9 M�  ۦ  զ  0y N	�   &�  $�  0w O	�   K�  I�   1 : =               �#  2�< =�  U2y: =+�  T2C: ==�   Q 3G          @      �Q  )Y  p�  n�  )e  ��  ��  )q  �  �  )}  =�  7�  4�  4�  4�  5G   	  )Y  ��  ��  )e  ��  ��  )q  ��  ��  )}  ٨  ר  * 	  +�  �  ��  +�  +�  %�  +�  v�  t�  #        E    $Ur $Ts  #        E     $Uz  #        �  D  $Uz $Qq $Rr  #        E  b  $Uz $Tt  #        �  �  $Uz $Tt $Qq $Rr  #        E  �  $Uz  #        E  �  $Uz  #        �  �  $Uz $Qq  #        E  �  $Uz $Tt  #        �  "  $Uz $Tt $Qq $Rr  #        E  :  $Ur  %        E  $Ur     3�
          �      �  )�
  ��  ��  )
  Ū  ��  )  �  �  )"  i�  c�  4.  4;  4H  5�
  p	  )�
  ��  ��  )
  ��  ��  )  ݫ  ۫  )"  �  �  *p	  +.  B�  *�  +;  B�  <�  +H  ��  ��  #        �  6  $Ur $Ts  #        �  N  $Uz  #        �  f  $Uz  #        T  �  $Uz $Tt $Qs $Rr  #        �  �  $Uz  #        �  �  $Uz  #        �  �  $Uz  #        T  �  $Uz $Qq $Rr  #        �    $Uz $Tt  #        �  2  $Uz  #        T  V  $Uz $Tt $Qq  #        �  n  $Uz  #        �  �  $Uz  #        �  �  $Uz  #        T  �  $Uz $Qq $Rr  #        �  �  $Ur $Tt  #        �  �  $Ur  %        �  $Ur     3�	          �      �]   )�	  ��  ��  )�	  ܭ  ֭  )�	  .�  (�  )�	  ��  z�  4�	  4�	  4�	  5�	  �	  )�	  ή  ̮  )�	  ή  ̮  )�	  ��  �  )�	  �  �  *�	  +�	  [�  A�  +�	  n�  h�  +�	  ��  ��  #        �
  �  $Ur $Ts  #        �
    $Uz  #        �
  $  $Uz  #        �
  <  $Uz  #        �	  f  $Uz $Tt $Qs $Rr  #        �
  ~  $Uz  #        �
  �  $Uz  #        �
  �  $Uz  #        �
  �  $Uz  #        �	  �  $Uz $Tt $Qq $Rr  #        �
    $Uz  #        �
     $Uz  #        �
  8  $Uz  #        �
  P  $Uz  #        �	  n  $Uz $Qq  #        �
  �  $Uz $Tt  #        �
  �  $Uz  #        �
  �  $Uz  #        �
  �  $Uz  #        �	  �  $Uz $Qq $Rr  #        �
     $Ur $Tt  #        �
  .   $Ur  #        �
  F   $Ur  %        �
  $Ur     37          �       �b!  )I  ߰  ݰ  )U  �  �  )a  Z�  T�  )m  ��  ��  4y  4�  4�  57  
  )I  ��  ��  )U  ��  ��  )a   �  �  )m  H�  F�  *
  +y  s�  m�  +�  ��  ��  +�  �  �  6�  P
  6	)�  �  
�  )�  e�  [�  *P
  +�  ܳ  س       3�          <      ��"  )�  �  �  )�  F�  @�  )�  ��  ��  )�  �  �  4�  4�  4�  5�  �
  )�  8�  6�  )�  8�  6�  )�  ^�  \�  )�  ��  ��  *�
  +�  ��  ��  +�  ��  ��  +�  $�  "�  7�          �
  �	)  N�  H�  )�  ��  ��  *�
  +  �  ��  +   k�  g�  ++  ��  ��       3�                 ��#  )�  ��  ��  )�  ׸  Ѹ  )�  )�  #�  )�  {�  u�  4  4  4  5�  0  )�  ɹ  ǹ  )�  ɹ  ǹ  )�  �  �  )�  �  �  *0  +  B�  <�  +  ��  ��  +  ��  ��  7*          �  �	)E  �  ٺ  )8  O�  ?�  *�  +R  4�  $�  +_  �  	�  +l  �  �  +w  4�  .�       3�          @      �%  )  ��  ��  )  ��  ��  )  �  
�  )*  b�  \�  46  4C  4P  5�    )  ��  ��  )  ��  ��  )  ֿ  Կ  )*  ��  ��  *  +6  )�  #�  +C  w�  u�  +P  ��  ��  7\          �  [	)w  ��  ��  )j  �  �  *�  +�  {�  w�  +�  ��  ��  +�  ��  ��  +�  �  �  +�  f�  ^�       3                �P&  )+  ��  ��  )7  ��  ��  )C  C�  =�  )O  ��  ��  4[  4h  4u  5     )+  ��  ��  )7  ��  ��  )C  	�  �  )O  1�  /�  *   +[  \�  V�  +h  ��  ��  +u  ��  ��  7�          p  �	)�  ��  ��  )�  v�  h�  *p  +�  C�  ?�  +�  }�  {�  +�  ��  ��  +�  ��  |�  +�  a�  S�  +�  8�  *�       3�          �       ��'  )�  �  �  )�  ,�  &�  )�  ~�  x�  )�  ��  ��  4�  4�  4�  5�  �  )�  �  �  )�  �  �  )�  D�  B�  )�  l�  j�  *�  +�  ��  ��  +�  ��  ��  +�  F�  D�  #        
  A'  $Uz $Tv $Qq $Rr  #        
  k'  $Uz $Tt $Qq $Rr  #        
  �'  $Uz $Tt  %        
  $Uz $Tt $Qq $Rr     3�          r       ��(  )�  r�  j�  5�  0  )�  ��  ��  #        +  (  $U	         "        +  #        �  9(  $Us $TD #        +  X(  $U	         "        +  #        �  �(  $Us $T( 8        +  $U	           3z          F       �E)  )�  +�  #�  5z  `  )�  ��  ��  #        +  �(  $U	         "        +  #        �  ()  $Us $T2 8        +  $U	           3�          �       ��*  )�  ��  ��  )�  �  �  )�  Y�  S�  )		  ��  ��  4	  4"	  4/	  5�  �  )�  ��  ��  )�  ��  ��  )�  �  �  )		  G�  E�  *�  +	  r�  l�  +"	  ��  ��  +/	  ,�  "�  #        ;	  **  $Ur $Tx  #        ;	  H*  $Ur $Tx  #        ;	  f*  $Ur $Tx  #        ;	  �*  $Ur $Tx  #        ;	  �*  $Ur $Tx  #        ;	  �*  $Ur $Tx  %        %+  $U	            9� � 	7	:    
 9� � 	69��  ��  d9�= �= Z9    9� � ! �   Q8  S#  :@ �*  ,�@     9      ��  O  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  9�  0t  4  e2    �0  }  ��  (  
K   J�  D   �C  
D  ���� �C  N\  ڵ  RP  ) �  J @4  � "�    � '
4  �� *	�   
 -D  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 �   D  =    �  
K   Y�  �?  N> �> i? �? ~? �? D@ A �? 	�@ 
 �@ eJ  Xi	@  �> m@   �> n	�   � sU  �� w\  �@ {q   c� \  (�@ ��  0�? ��  89> ��  @? ��  Hs> ��  P �  �  U  �   F  [  �   q  D   b  �  �   �   �    w  �   �  D  �   �   �    �  �  �    �  �  �  �    �  �  D  �    �  u@ ��  h�	�  �> �@   �> �	�   � ��  �� �\  d> ��   C> �\  (Z@ �\  0�? ��  80? ��  @%? ��  H�> �\  P�> ��  X�@ �\  ` �  �  R   �  R   �    �  �  R    �  �  R   �   �  f@ ��  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   �  	��  ��   	�\  ��  	�  �{  �  	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  �Q  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   	�  	�   	q  	*  �   	��  
%�   !  '	�7e     -  ,	�7e     9  1	�7e     E  5	�7e     �@ 9�  	��e     �  �> :�  	��e     �    <	�7e     	  =	�7e     	> B�  	�@ C�  	�@ D�  	�= E�  	@ I�   	�> M�   �  8  =     �@ \(  �  T  =     �? gD   ��> �	�  R�@            ��> �B�@            �#? �2�@            �  t �R   ��  ��  ? �'�  �  �  A�@     U�UT�T  .? �"�@            �K  t �R   _�  Y�  1�@     U�U  �? �R   �@            ��  "8 �R   ��  ��   len �&�   �  ��  �@     U�UT�T  �? ~ �@            �M? v��@            �b> n��@            �-	  Ml  n�   U�  O�  �@     U�U  Y? i!�	 e�= ]Ƈ@            ��	  �> ]"D  ��  ��  �> ].�   ��  ��  ݇@     U�UT�T  
? Q	�  ��@            ��	  v? Q�   K�  E�  Ç@     U�U  7> I��@            �2
  v? I�   ��  ��  ��@     U�U  �? <�   f�@     >       �6  �@ <D  ��  ��  v? <*�   A�  ;�   vol <7�   ��  ��   sep <@�   0�  (�  ��@     U�UT�TQ5�Q�Q $�O$,( 0�Q�Q $�O$,(  $0*( R7�R��R $� $,( 0�R��R $� $,(  $0*(   �@ 31�@     5       �  v? 3�   ��  ��   vol 3+�   �  �   sep 34�   ��  ��  e�@     U�UT5�T�T $�O$,( 0�T�T $�O$,(  $0*( Q7�Q��Q $� $,( 0�Q��Q $� $,(  $0*(   "> C  #vol (C  #sep 2C   �   ?? �@     B       ��@ �   ݆@            ��  �@  D  S�  M�  �@     U�U  $@ ���@     8       �%� �,�@     y       �8  &�> ��  ��  ��  '"@ ��  ��  ��  '�> ��  .�  *�  '/> ��  ~�  x�  (P  ��@     ��@            ��  )]  ��  ��  *��@            +i  �  �    (8  ��@     ��@            ��  *��@            +E  5�  3�    ,:�@     �  �  U	�B      ,G�@     �    U	&�B      ,S�@     �  *  U	-�B      -|�@     �   .*@ �P  /i �	�    .> �t  0�> �#�  /i �	�    1�= r�  �  0< r,�  0*  rA@  2len s$�   /i u	�    36	  އ@            �4� � 	!4�C  �C  A G   �;  S#  PE �*  e�@           {�  �P  �)  �=   ,	  int ^&  9�  nC (g   �E p   �   �   =     	D  �   
�E  �    
�G  �   
F  K   
3E  K    �  �1  @G  Q  G   �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2D   8;:  5D   < M  1  �K 8"�   �  Kl  T  �  Ll  �  Ml  *  c[   0t  �  e2  �    �0  }  C ��  G  8J �G  �D �D   �G �D   7G �D   ��  �  �   	J5  D   �C  
D  ���� �C  	N  ڵ  	R  �  
D   q  
�  ��  %G  q  : �D   3 �D   � �D   � �D   O �D   �
 �G  A  ��  �G  �\  �5  �  ��  �  ��  �D   ��  �D   2�  �5  ��  �D   Ɇ  ��  ��  �D   ��  �D   �h  �D   rK  �D   l�  �D   ]�  �D   ��  �D   w
 r  =� �  ��  .�  ^�  2[   }�  7�  �� ;�    	�  r�     .� $%  O� )I       G   �  �  %       1   I    �   K   1    +  ��  ,�  O  oS  'm  dS  ()�  � +
�   � ,  @�  -
D   >z .
D   �  /K   �H  3�    M  �  =    a  �� 7�  �� 8�   �F >#  �F @8  ڈ B�   �C C5  �H  D8   �  �D G8  	��e     G e5  	��e     �  {  =   	 k  �G �{  	h�B     B �{  	X�B     �E �{  	H�B     �  �  =   	 >G ��  	��e     �B �  	 8e     �  �H �	5  �@     �      �t  82  �'�   _�  Y�  �| �5K   ��  ��  >z �@D   �  ��  �� �5  	�7e     �@     �       p �D   P�  L�  i �D   ��  ��  val �D   ��(�@     t  �   U	+�B      T1 X�@     �     U  T	3�B      t�@     �  8   U  T	:�B      ��@     �  ]   U  T	@�B      !،@     �   T��   "��  g?�@     8      ��
   gG  ��  ��  #�F i
�
  ��zJ j�  ��z$#G k8  ?�  =�  $�C l5  d�  b�  %�
  ��@     ��@     �       �	�	  &�
  ��  ��  ��@     �       '�
  (�
  ��  ��  (�
  ��  ��  %1  ��@     ��@     
       J
�  !Ê@     �   U	��B       %�
  ˊ@     ˊ@     X       O;	  &   F�  B�  ˊ@     X       (  ��  �  (  ��  ��  (%  h�  b�  )�@     �  !�@     �   U	��B      Ts 8$8&   @�@     �  S	   Us  ]�@     �  �	   U|  Ts  Q	��B      R	��B      Xv  e�@     �  �	   U|  m�@     �  �	   U|  !u�@     �   Uv    Չ@     �  �	   U	L�B      $�@     �  
   Tv  Q��z 5�@     �  4
   U	z�B      )A�@     �  ��@     �  m
   U|  T
  Qv  R��z !��@        U	}�B       M  �
  *=   � +A CD   �
  ,|G C!G  -��  E	D   -tG FG  -&E GG  -GA H1    +�J G  1  ,b[ &G  -��  G  .r G  .s G   /�C D   0/ �(�@            �r  1#G �8  ��  ��   2aH �	5  3� ���@     -       �  4�_  �!G  ��  ��  )�@       �@     m  �   U�h )�@       �@          U	6�B      5%�@        3	 �و@            �m  6i �	D   �  �  �@       Y   U= 7��@        U:  3H ���@     E       ��  8msg �G  ��  ��  6i �	D   ��  ��  1�A �	D   ��  ��  ˈ@       �   U  7و@     &   U�U  9�C ��  w�@     u       �_  4>z �_  (�  "�  1B ��  |�  t�  :^J �	D   1qH �D   ��  ��  6p �	D   ��  ��  ;e  ��@     ��@     '       �  <�  <�  &v  $�  "�  ��@     '       (�  O�  G�  ��@     �  �   U
s D$ $ & !ҋ@     t   U	ٕB      Ts   ��@     t  0   U	ՕB      T1 )��@     2  !�@     >   U	�B      T|   D   =?F _�  �  >>z _#_  >qH _-D   >^J _>D   :B a�   3�D W��@            ��  ?on WD   U?off WD   T@9F W%D   Q 3 Ie�@     .       �]  4ڈ I�  ��  ��  4�C I+5  �  ��  1#G K8  O�  M�  !w�@     �   UH  Ar  %�@            �B��  ��  
%B:�  :�  BSJ SJ "	BC C OB��  ��  ABZH ZH #BG�  G�  /Bm�  m�  @C�E �E  B�J �J iB�= �= ZB�F �F .B?J ?J 
+	C     B� � ~B    B� � (B��  ��  d 6   �?  S#  �K �*  }�@     X       ��  �U  ,	  e2    �J R   �  �0  }  int ^&  K F   UK 
�   u   K "u   	��e     R Yԍ@            �	sK SӍ@            ��   
r� Sg   U 	B�  K΍@            �7  ms Kg   v�  r�  Ӎ@     !  U�U  @ =g   ��@            ��  G ?u   ��  ��  �  ��@        A��@     -     *g   ��@     +       ��  G ,u   ��  ��  �  ��@     �  .��@     -    �K %g   �  }�@            �!  ��@     -   JK JK }K }K 
 8   A  S#  �K �*          �      '�  W  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  9�  �K 4  �K   �  
buf !   L "	1   Q #	1   @�  $K   /  %   K   �  �K  �K L  �K �  K   "�  ��  WH  �~  �O  �m  ��   �  ��  ��  	 K     �K   L  CL �  "  e2  RL ��           :       ��  
 ��  5�  1�  @�  �,D   v�  n�  <L �@�  ��  ��  �K �K   �  �            U	          (  lL �D                  ��  
 ��  U 1L �               �C  
 ��  W�  O�                      U�U  �K �               ��  
 ��  Ubuf �*�  TL �7�  Q R   1   �L k1           �       �n  ptr kn  ��  ��  >z k+1   �  �  +L k81   K�  E�  
 kH�  ��  ��  ��  m	1   ��  ��          .       �K {  B�  >�          $  _  T1Q0             t  \L Z
�          K       ��  � \�  ~�  x�          $  �  U T1Q0         $  U
 T1Q0  �K :1           Y       ��  buf :R   ��  ��  >z :$1   8�  .�  +L :11   ��  ��  
 :A�  4�  ,�  ^� <	1   ��  ��          0  U	          vL *
�          -       �  buf *R   ��  ��  L *+1   ;�  5�  � ,�  ��  ��          $  U T1Q0  ��  ��  d� � 7	� � 6      l   �B  S#  �L �*  Ս@     �       ��  �W  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"R   �  K  �   �  L  �  M  9�  e2    �0  }  	K   Jf  
D   
�C  
D  ���� �C  NB  �  �   q  �  �   r  	 Df     ~  		(Df     �L ��   5�@     &       �  sep ��   ��  ��  M�@     W  Us T/  �  �4�@            �/  i ��    �L KI  �L K"�    � D�    �@            ��  Wy D�   ��  ��  $�@     �  U�UT0  ?J ?	f  $�@            ��  Wy ?�   �  �  *�@     I  U�U  ��  +�   Ս@     K       �W  Wy +�   O�  I�  �L +*�   ��  ��  i -	�   ��  ��  �@     c  U~   ��  ��  &:�  :�   �    >D  S#  #M �*  [�@     =       f�  �Y  t�   =   int k   k   �L  M M �L  �  �L $v�@     "       ��   box %�   Ux &1   Ty '1   Q 	1   
�L [�@            �box �   U  �   �D  S#  9M �*  ��@     �       ��  �Y  �)  �=   ,	  e2    �  �0  }  int ^&  R   J�   D   �C  
D  ���� H#	�   	� '
�    	�^  (1    	.�  )	g   (	o�  -1   0	i�  .	g   8	��  /
  < 
    =    1  
    =    �  0�   ,M R'�@            �k  cht Sk  C�  =�  �< T
q  ��  ��       �~  #g   ��@     �       �cht $k  ��  ��  key %	  T     �E  S#  R �*  8�@     8      t�  �Z  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  �   	int �   �K 8"T   
�  K  �   
�  L  
�  M  9�  
uO 	�   
YP �   
kS �   e2    �0  }  K   J�  D   �C  
D  ���� �C  Nr  
�  �   
q  �  �   ��  -�   	0Df     GR 1�   	��e      U 2�   	��e     K   5/  ~M   P �T R eN  VN ;   =	�  � @�    ;Q CR   *� F/  �U K	�   �M Q	�   eS U�   OP V;  X	�  
T Z�   �T [	�   ��  \�    �  �P ]�  �  �  =   K �M o�  	@Ge     �T ��  	 Ge     �  /  =   v QS �  	@8e     T �  	 8e     �   m  =    ]  �Q 4m  	��B     N '�   ,�@     D       �S  �  '�   	�  �  �e  )�   H�  B�  B�@     
  �  U	|�B      Q�@         T	 �B     Q0 \�@     "  1  Us  k�@     .  U	*�B     Ts   � �@     J       �  dir �   ��  ��    �@     �@            �  �@              ��  ��  ��@     :  U2   �@     .  �  U	��B       ,�@     "   !�T ��   -  "��  ��    �R ��  ��@     $       ��  � � �   ��  ��  �R ��  2�  0�  đ@     �  U�U  �  #N ��  ��@     %       ��  � �$�   Y�  U�  �R ��  ��  ��  ��@     �  U�U  �   JU ��   v�@     #       �c  � ��   ��  ��  �R ��  ��  ��  |�@     �  U�U  �M �	�  �@     �       �  � ��   �  �  �| �)�   \�  V�  �R ��  ��  ��  #�
  ��@     0  �i  $�
  �  �  $�
  7�  1�  %0  �
  ��  ��  �@     
  #  Uv  /�@     �
  ;  Uv  ;�@     �
  S  Uv  a�@     F  Uv    �@     �  U�U  � �ː@            ��  � ��   ��  ��  ;Q �'R   �  �  �R ��  _�  ]�  Ԑ@     �  U�U  &N ��  ~�@     F       ��  � �+�   ��  ��  ��  ��  ��  ��  ��@     �
  e  U	 Ge     Tv  ��@     �
  �  U	 8e     Tv  ��@     R  U	r�B     Tv   � Y�@     �       ��	  'i [	�   j�  b�  �@     ^  	  U	��B     T1 C�@     .  !	  U	��B      \�@       8	  Q0 v�@     .  W	  U	��B      ��@     ^  {	  U	ǖB     T1 ��@     .  �	  U	ԖB      @       Q0  �T @�@            �
  (`R @$�   U( P @0�   T[R B�   ��  ��  P C�   ��  ��   )|Q 6� ,��@            �^
  (OR ,!�   U((U ,4�   T *�O �z
  +�U �9z
   �  *�M ��
  ,def �$�  +�| �/�   "tQ �	�    !�R ��   �
  +Q �$�   "��  �	�    *qP I�
  +�U I9z
   &�S �  8�@     F       �t  �U :z
  &�   �  � L�   x�  r�  'i 	�   ��  ��  j�@     j  U~   -�
  ď@     9       ��  $�
  �  �  .�
  �l/�
  ӏ@            �  $�
  ��  }�  ӏ@            .�
  �l  0�@     v   1
  �@            �2��  ��  	2��  ��  +2xT xT 2��  ��  d2��  ��  	A2�M �M 	'2��  ��  
72��  ��  %2'�  '�  2�Q �Q h *    I  S#  �U �*  p�@     J      ��  �^  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"R   �  K  �   �  L  �  M  e2    �0  }  ��  %�   	<]  �   	XRe     	��  �   	TRe     	h  �   	PRe     	��   �   	LRe     	�  !�   	HRe     	�j  "�   	DRe     	��  #�   	@Re     	v  $�   	<Re     	R  %�   	8Re     	��  &�   	4Re     	�U  ,�   	0Re     	�n  -�   	,Re     	�  .�   	(Re     	��  0�   	$Re     	�  1�   	 Re     	��  2�   	Re     	u  4�   	Re     	_b  5�   	Re     	N  6�   	Re     	�o  <�   	Re     	�T  >�   	Re     		�  ?�   	Re     	^�  @�   	 Re     	��  A�   	�Qe     	��  B�   	�Qe     	�  C�   	�Qe     	[n  D�   	�Qe     	��  E�   	�Qe     	�  P�   	�Qe     	��  Q�   	�Qe     	0h  R�   	�Qe     	�g  S�   	�Qe     	��  T�   	�Qe     	^�  U�   	�Qe     	�a  V�   	�Qe     	>�  W�   	�Qe     	��  X�   	�Qe     	��  _�   	��e     	��  `�   	�Qe     	�P  a�   	�Qe     	#L  c�   	�Qe     	gz  e�   	�Qe     	�  f�   	�Qe     	�k  g�   	�Qe     	�  h�   	�Qe     	Ӄ  j�   	�Qe     	�v  k�   	�Qe     	O  n�   	�Qe     	��  o�   	�Qe     	-�  p�   	�Qe     	��  q�   	�Qe     	Ϊ  u�   	�Qe     
�   �  =    	��  v�  	@Df     	ӄ  z�   	�Qe     	r�  {�   	�Qe     	~�  |�   	�Qe     	��  }�   	�Qe     	��  ~�   	|Qe     	��  �   	xQe     	��  ��   	tQe     	��  ��   	pQe     	��  ��   	��e     	J�  ��   	��e     	Ei  ��   	lQe     	��  ��   	hQe     	��  ��   	dQe     	A�  ��   	`Qe     	��  ��   	\Qe     	��  ��   	XQe     	��  ��   	TQe     	 t  ��   	PQe     	��  ��   	LQe     	!�  ��   	HQe     	oa  ��   	DQe     	/z  ��   	@Qe     	��  ��   	<Qe     	1P  ��   	8Qe     	�  ��   	4Qe     	Ʒ  ��   	0Qe     	�T  ��   	,Qe     	�o  ��   	(Qe     	�b  ��   	$Qe     	~�  ��   	 Qe     	��  ��   	Qe     	�S  ��   	Qe     	��  ��   	Qe     	U  ��   	Qe     	Dl  ��   	Qe     	��  ��   	Qe     	��  ��   	Qe     	�p  ��   	 Qe     	"�  ��   	�Pe     	�  ��   	�Pe     	�K  ��   	�Pe     	��  ��   	�Pe     	�  ��   	�Pe     	tW  ��   	�Pe     	'�  ��   	��e     	�a  ��   	��e     	�W  ��   	�Pe     	̶  ��   	�Pe     	�`  ��   	�Pe     	��  ��   	�Pe     	��  ��   	�Pe     	̨  ��   	�Pe     	��  ��   	�Pe     	�X  ��   	�Pe     	��  ��   	�Pe     	��  ��   	�Pe     � ���@            � wh�@     Q       ��  �  w&K   ��  ��  � y
�  �@i zK   �  �  ��@        S  U	��B     T	�Qe      ��@     !   �  Uw T Q	��B     Rs ��@        Uw Ts2$@Df     "  
�   �  =    # X�@     y      �#  ��@          U	W�B     T	<Qe      �@        2  U	i�B     T	8Qe      �@        ^  U	u�B     T	4Qe      ,�@        �  U	��B     T	0Qe      ;�@        �  U	��B     T	,Qe      J�@        �  U	��B     T	(Qe      Y�@          U	��B     T	$Qe      h�@        :  U	��B     T	 Qe      w�@        f  U	КB     T	Qe      ��@        �  U	ߚB     T	Qe      ��@        �  U	�B     T	Qe      ��@        �  U	��B     T	Qe      ��@          U		�B     T	Qe      @        B  U	�B     T	Qe      ј@        n  U	)�B     T	Qe      ��@        �  U	8�B     T	 Qe      �@        �  U	I�B     T	�Pe      ��@        �  U	[�B     T	�Pe      �@          U	j�B     T	�Pe      �@        J  U	x�B     T	�Pe      +�@        v  U	��B     T	�Pe      :�@        �  U	��B     T	�Pe      I�@        �  U	��B     T	��e      X�@        �  U	��B     T	�Qe      h�@        U	��B     T	�Qe        H9�@     �       �O  I�@        n  U	؛B     T	lQe      X�@        �  U	�B     T	hQe      g�@        �  U	��B     T	dQe      v�@        �  U	�B     T	`Qe      ��@          U	�B     T	\Qe      ��@        J  U	�B     T	XQe      ��@        v  U	ɛB     T	TQe      ��@        �  U	-�B     T	PQe      ��@        �  U	=�B     T	LQe      З@        �  U	L�B     T	HQe      ߗ@        &  U	Y�B     T	DQe      �@        U	f�B     T	@Qe       g 3e�@     �       ��  u�@        �  U	x�B     T	�Qe      ��@        �  U	��B     T	�Qe      ��@        �  U	��B     T	�Qe      ��@          U	��B     T	�Qe      ��@        J  U	��B     T	|Qe      ��@        v  U	��B     T	xQe      ϖ@        �  U	��B     T	tQe      ޖ@        �  U	̜B     T	pQe      �@        �  U	؜B     T	��e      ��@        &  U	�B     T	��e      �@        R  U	��B     T	�Pe      �@        ~  U	ΙB     T	�Pe      )�@        �  U	�B     T	�Qe      9�@        U	0�B     T	�Qe       �U 7�@     .      ��  ��@          U	ɞB     T	Re      ��@        J  U	��B     T	$Re      ��@        v  U	ǟB     T	 Re      ��@        �  U	|�B     T	Re      ��@        �  U	��B     T	Re      Ε@        �  U	��B     T	�Qe      ݕ@        &  U	�B     T	�Qe      �@        R  U	*�B     T	�Qe      ��@        ~  U	6�B     T	�Qe      
�@        �  U	A�B     T	�Qe      �@        �  U	L�B     T	�Qe      (�@          U	X�B     T	�Qe      7�@        .  U	��B     T	�Qe      F�@        Z  U	��B     T	�Qe      U�@        �  U	-�B     T	�Qe      e�@        U	c�B     T	�Pe       V  ��@     �       ��  ��@        �  U	ɞB     T	Re      ��@        &  U	-�B     T	�Qe      ��@        R  U	c�B     T	�Pe      ͔@        ~  U	��B     T	Re      ܔ@        �  U	�B     T	Re      �@        �  U	�B     T	 Re      ��@          U	&�B     T	�Qe      	�@        .  U	;�B     T	�Qe      �@        Z  U	M�B     T	�Qe      '�@        �  U	d�B     T	�Qe      7�@        U	q�B     T	�Qe       V ��@     �       �V  �@        �  U	ҞB     T	0Re      &�@        %  U	ܞB     T	,Re      5�@        Q  U	�B     T	(Re      D�@        }  U	��B     T	$Re      S�@        �  U	�B     T	 Re      b�@        �  U	�B     T	Re      q�@          U	c�B     T	Re      ��@        -  U	o�B     T	Re      ��@        U	��B     T	Re       C
 �p�@     �      �   ��@        �  U	y�B     T	XRe      ��@        �  U	��B     T	TRe      ��@        �  U	��B     T	PRe      ��@        $  U	��B     T	LRe      ��@        P  U	��B     T	HRe      ˒@        |  U	��B     T	DRe      ڒ@        �  U	ԟB     T	@Re      �@        �  U	ݟB     T	<Re      ��@           U	�B     T	8Re      �@        ,  U	�B     T	4Re      �@        X  U	�B     T	��e      %�@        �  U	�B     T	�Qe      4�@        �  U	�B     T	�Qe      C�@        �  U	9�B     T	��e      R�@          U	C�B     T	�Pe      a�@        4  U	O�B     T	�Pe      p�@        `  U	X�B     T	�Pe      �@        �  U	��B     T	�Pe      ��@        �  U	��B     T	�Pe      ��@        �  U	��B     T	�Pe      ��@          U	ޙB     T	�Qe      ��@        <  U	�B     T	�Qe      ʓ@        h  U	�B     T	�Qe      ٓ@        �  U	�B     T	�Qe      �@        �  U	B�B     T	�Pe      ��@        �  U	M�B     T	�Qe      �@        U	��B     T	�Qe       � � G�  G�  / 5   rJ  S#  @V �*  ��@     L       ��  �_  ,	  int ^&  9�  e2    �  �0  }  2V ?   k� p   t�   8   H_  /	�   ̙@     :       ��   a /�   Ub /%�   I�  E�  ��@            	��  7
|   ��  ��    
d  "�   ��@            �a #�   ��  ��  b $�   T  *z   *K  S#  �[ �*  p          ��  �`  �)  �9   ,	  int ^&  9�  �  �1  @�   Q  �    �   	-   62  #	-     &	-   �5  )	-    �@  ,	-   (.  -	-   0*  2@   8;:  5@   < �   1  �K 8"^   	�  K  �   	�  L  	�  M  0t  0  e2    �0  }  ��  $  
W   J|  D   �C  
D  ���� �C  NX  ڵ  RL  �  
W   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
W   /  ��   [r  �4 #�  �   �X  5�  
W   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K)  
@   P�  =_  ��   R�  N�  ��  ��   �p  W�  
W   3�  ��   ({  ��  ğ   F]  8�  
W   ;U  �  � | 7	  �
 ` � � � 	 � F
  
W   Y�  ��   �c  |  ��  l  ��  �   
W   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {�  
W   �*  &�   �  º  GY  �f  ��   v�  ��  
W   �o  GQ   ϼ  �  �_  X  &�  �b   �   z   	Y�  	%o  	��  	&o  	� 
.U  	"|  *|  	��  +|  	I�  ,|  	�a  -|   	Z  ��  ">   E�  #>  e% $E  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	@   a  2
�  �T  3
�   Mx 4�  
W   !�  �p   �  ��  S�  ��   �F  'f  *	�  *� ,�   "G  C	@   (G  C@   �]  C@   :G  C@    �U  D�  �  �  	��  ��   	�\  �|  	�  �'  �  	��  �@   	��  �@   	2�  �|  	��  �@   	Ɇ  ��  	��  �@   	��  �@   	�h  �@   	rK  �@   	l�  �@   	]�  �@   	��  �@   (		  ��  E      E  Vd  !E  �  "E  �� #	   @     9    � %�  @   5  9    	N�  %%  	��  '�    =� _  ��  .�  ^�  2!   }�  7�  �� ;W    	�  r�  �   .� $�  O� )   �  �  �    S  �  �  �   �  -     �  W   G   -    �  ��  ,�    oS  '3  dS  ()�  � +
�   � ,�  @�  -
@   >z .
@   �  /G   �H  3�    �   �  9    '  	�� 7�  	�� 8W   
W   "	  ��  WH  �~  �O  �m  ��   �  ��  ��  	 t�   @   	  	  $	  9   �' 	  	��  1$	  	]  4A	  	  	  X	  9   � G	  	Zy  8X	  �  	  9   9   � i	  	��  ;	  Ʃ  QW   �	  �	  �	  9     �	  	�  W�	  �p  #�	  �	  �	   S�  $�	  �	  �	  G    T}  %
  
  
  G   G    '	I
  acv )�	  ��  *�	  ��  +�	   �y -
  �Y  6I
  ��  :�
  s�  <�
   �H  =�
  xz  >U
   a
  x @a
  E  �
  9    7  �
  9    
�	  x �E   y �E  Mp �E  *� �E  ޽  �E   ~x ��
  
W   l  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �  
W   ��'  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  ux   (x	y(  !�u zl   !� {	@   !s |	@   !� ~I
  !N�  �'  !��  �	@   !��  �	@     J]  �(  y(  �(  9   � "�^  ��(  "�  �o  #W   ��+  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �(   \	W-  !�Y  	@    !*O  	@   !��  	@   !�  	@   !b�  	@   !��  	@   !�  	@   !+�  	@   !Zp  	@    !o�   	@   $!m�  !	@   (!4�  "	@   ,!�  #	@   0!�  $	@   4!��  %	@   8!L� &	@   <!��  '	@   @!  (	@   D!��  )	@   H!\q *	@   L!z�  +	@   P!�  ,	@   T!/�  -	@   X ʤ  /
,  W-  t-  9   � "��  1d-  �]  ��W/  `e ��
   x �	  y �	  z �	   ��  �W/  (cN  �W/  0Mp ��	  8�u �l  <� �@   @�H  �W/  Hr�  �W/  P��  ��/  X��  �	  `m�  �	  d��  �	  h  �	  l3F  �	  p8F  �	  t=F  �	  x��  �@   |*� ��+  �y� ��/  �s �@   ��� ��/  ��  �@   ��  �@   �ʺ  �@   ��l  �@   �! �  W/  �!��  @   �!��  	@   �!�R  ~1  �!f�  @   �!I}    �!��  W/  � �-  Gx  ��/  >} �4   �}  �E  �|  �E  
 ]/  W-  y(  $d  HN~1  mo P�2   ��  Q�9  cmd RZ  �  W	  (_  Y	   #_  [	  $bob ]	  (�  a@   ,�[  b@   0sb  d@   4d]  g�9  8�W  h�9  P��  i|  h�� l%  l�N  m�  |E�  p�  ��W  r�9  �~�  s%  �*� t%  ��� w@   ���  x@   �X�  |@   ��e  @   ���  �@   �g  �@   ��u  �@   �|G ��   �Q  �@   ��  �@   �o�  ��2  �%�R  �@    %��  �@   %�  �@   %h  �:  %I�  �|  @ �/  �z �-  C	�1  x E	   y F	   �{ H�1  (T	�1  `e V�
   x W	  y X	  z Y	    	�  [�1  �a	�2  = c	   F�  d	  �~ eE  h�  fE  
t�  gE  �k hE  tag iE  �N  l
@   ��  o�2  ��  r
%   iK  u�1  0��  x
@   XS�  {�2  `��  ~G   h��  �@   pu| ��3  x �1  �}  X��3  v1 �V4   v2 �V4  dx �	  dy �	  �  �E  �k �E  tag �E  �W  ��
  �o �\4  $��  �J4  4SX  �4  8d�  �4  @��  �
@   H��  �G   P �3  �2  �z �2  �	4  2�  �	   ]  �	  �h  �E  �N  �E  
�K  �E  >} �4   �3  �}  ��3  
W   �J4  ��   �  o�  ��   ��  �#4  �1  	  l4  9    �u  ��2  �z �]/  8�	�4  v1 �V4   v2 �V4  82  �	  Mp ��	  [�  ��4   �  ��4   SX  �4  (d�  �4  0 4  l4  A{ ��4   4	e5  &x 	   &y 		  &dx 
	  &dy 	  !�o e5  !)�  �
  0 	  {5  9   9    (} 5  �  *�  'v  @2J6  !@�  4J6   &x1 5@   &x2 6@   !.]  8	  !5]  9	  !�� :	  !��  =@   !�  @	   !��  C	  $!�n  GP6  (!9x  HP6  0!�^  IP6  8  5  E  >�  K�5  '�h  PR?7  !s�  U?7   !�H  V?7  &x1 X@   &x2 Y@   &gx \	  &gy ]	  &gz `	   &gzt a	  $!�x  d	  (!� f	  ,!~�  i	  0!t  k	  4!.� l@   8!�  pE7  @!	�  r@   H c6  �5  �h  tc6   �	�7  !�c  �|   !�O  ��7  !�x  �
�7   E  �7  9    �  �7  9    I�  �X7   �	�7  !�  �@    !�  ��7   �7  �  ��7  (��	�8  !  �	   !�  �	@   !t�  �	@   !��  �	@   !/�  �	@   !�  �	�  &top �	�8  )��  �	�  U)��  �	�  V)� �	�8  W)�  �	�  � �  �8  9   ? ��  ��7  	9  ~�  *   �S  
@   ��   
@     !
@   �g  "
@   �^  #
@    ��  %�8  9  09  9    	S�  ' 9  
W   7]9  {�   U�  ~�   >	�9  �� @�/   s A
@   sx B	  sy C	   Nz E]9  
W   1�9  ��   ��  ��   �y  9�9  @   �9  9    |  �9  9    |  :  9    �9  :  9    hy ��/  (�	�:  in �|   d  �
@   �x  �
@   D  �
@   5O  �
@   �� �
%  �a  �
@   $ ��  �:  ��	';  2�  �
@    I�  �|  r�  �
@   �H  �
@   *F  �
@   ��  �
@   	�  �
@   ѵ  �
@   ��  �
@    F� �
@   $�  �';  ( �:  7;  9    ޴  ��:  	.L  &O;  	  	׮  )O;  	�  +O;  	�  ,O;  	�Q  .E7  	��  0@   	��  1@   	(_  2@   	դ  4@   	�j  7�;  @   	��  8�;  	@�  <@   	�O  =@   	(g  >@   	�^  E@   	�u F<  �7  	��  H@   	��  IV4  	��  K@   	a� LJ6  	w�  N@   	P{ O4  	��  Q@   	��  Ru<  x4  	��  T@   	�� U�<  {5  	�}  W@   	u| X�4  	M�  Z@   	P�  [�4  	��  a	  	��  b	  	�  c	  	�p  e�	  	�T  f=  :  	�a  j�	  @   (=  9   � 	ը  l=  �	  E=  9   @ 	�p  m4=  	 �  p	  	p|  q�	  	$Y  v@   	�K  y@   	g  {�=  �8  	d�  |�=  	��   	  		�  !	  	�3 #@   	_  $@   	-�  (@   	�f  )@   	�G  +	  	`�  ,	  	A�  -	  	��  /@   	��  1@   	P�  2@   E7  E>  9   9   / 	��  E/>  E7  a>  9   / 	Ԁ  FQ>  E7  �>  9   9    	7� Gm>  	�R  I@   	��  JE7  	��  U@   	P�  \�  	��  ]�  	L�  ^�  	ߵ  _�  	�  a�  	@�   J6  	[�   �4  	 �   �4  	SX   4  	d�   4  	��   @   	_�    @   	��   "|  	��   %|  	'�   &|  	�]   (|  V6  �?  9   � 	�P   *s?  	ӯ   +�?  V6  	|   -�?  E7  	��   .�?  	��   /�?  �?  �?  @   @    	��  !P6  �  ! �?  	qY  !"�?  	�  !#�?  E  "@  9   ? 	��  !%@  	��  !&@  	  J@  9   � 	@Y  !(:@  	  g@  9   ? 	V�  !)V@  K7  �@  9    	�h  "s@  	�  "�@  K7  	�  "K7  	�f  "!@  	r�  ""@  	��  "%P6  	��  "&P6  	׆  "'	  	��  "(	  	�  "*	  	��  "+	  	�  #E7  	��  #@   	�_  #@   	�_  #@   	b  #	  	t  #	  	j�  #"�  	�  #:@   	��  #;@   	��  #<@   	�W  #>E7  	hn  #@	  	U~  #A	  	�  #B	  	 �  #C	  	%�  #F�  	�u  #H�  	z  #I�  �   �A  9   	 	~ $8�A  	� %M@   	5 %N@   	�  &@   	q  &1B  �   	<]  '@   	��  '@   	h  '@   	��  '@   	�  '@   	�j  '@   	��  '@   	v  '@   	R  '@   	��  '@   	�o  ' @   	�U  '"@   	�n  '#@   	�  '$@   	��  '%@   	�  '&@   	��  ''@   	u  '(@   	_b  ')@   	N  '*@   	�  '-@   	��  '.@   	0h  '/@   	�g  '0@   	��  '1@   	^�  '2@   	�a  '3@   	>�  '4@   	��  '5@   	O  '7@   	��  '8@   	Ϊ  ':@   	��  ';	  	ӄ  '=@   	r�  '>@   	~�  '?@   	��  '@@   	��  'A@   	��  'B@   	��  'C@   	��  'D@   	�T  'F@   		�  'G@   	^�  'H@   	��  'I@   	��  'J@   	�  'K@   	[n  'L@   	��  'M@   	-�  'O@   	��  'P@   	��  'Q@   	J�  'R@   	Ei  'T@   	��  'U@   	��  'V@   	A�  'W@   	��  'X@   	��  'Y@   	��  'Z@   	 t  '[@   	��  '\@   	!�  ']@   	oa  '^@   	/z  '_@   	��  'c@   	1P  'd@   	�  'e@   	Ʒ  'f@   	�T  'g@   	�o  'h@   	�b  'i@   	~�  'j@   	��  'k@   	�S  'm@   	��  'n@   	U  'o@   	Dl  'p@   	��  'q@   	��  'r@   	�p  's@   	"�  't@   	�  'u@   	�K  'v@   	��  'w@   	�  'y@   	tW  'z@   	'�  '{@   	��  '}@   	��  '~@   	�P  '@   	#L  '�@   	gz  '�@   	�  '�@   	�k  '�@   	�  '�@   	Ӄ  '�@   	�v  '�@   	�a  '�@   	�W  '�@   	̶  '�@   	�`  '�@   	̨  '�@   	��  '�@   	��  '�@   	��  '�@   	�X  '�@   	��  '�@   	��  '�@   	
 (:  	 (;|  ) )wG  J @)H  � )"�    � )'
H  �� )*	@   
 )-H  �9 )0	@    Ml  )3	@   $	
 )8	@   (C� );	@   ,� )?	@   0� )BG   8 �   H  9    kG   )H	[H  � )K�    C� )N	@   "8 )QG   t )TG    . )VH  rH  @    gH  	: )�@   	3 )�@   	� )�@   	� )�@   	O )�@   	�
 )��   kG  �H   	R *�H  [H  �H   	� *�H  
W   *r�K  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	 +V@   Z  	��  ,M|  	(h  ,N@   	l�  ,N@   	�  -.|  	�  -/|  	�  -0|  	�  -2|  	w�  -8  	�  -9�  	�  -:�  	�_  -;�   	��  ->|  	�  -J|  	"�  -R�  	t�  -S@   	�w  -T@   	؜  -Y@   	q�  -[|  	Ƚ  -^�  	�  -_@   	�y  -`@   	b�  -c@   	+�  -f|  	��  -i|  	֘ -l@   	�J  -x@   	��  -y@   	ks  -@   	�  -�@   	J�  -�@   	�i  -�@   	��  -�|  	��  -�|  	��  -�|  	<� -�|  	��  -�|  	��  -�|  	5�  -�|  	<m  -�@   	 K  -�@   	�R  -�@   	op  -�@   	�m  -�@   	D  -�@   	X�  -�@   	If  -�@   	� -�@   	��  -�|  	�U  -�|  	`  -�|  	J�  -�|  	��  -�|  	� -��  :  /N  9    	�  -�N  |  KN  9    	� -�;N    gN  9   	 	,�  -�WN  	R�  -�N      �N  9    	�u  -��N  	��  -�7;  	�e  -��   �   �N  9   � 	(�  -��N  	�  -�|  "��  -�  "�v  -@   "n�  -@   "4�  -@   "*b -@   "��  -�K  	B .8@   	x	 .9@   M  XO  9   > 	D >HO  	�5 ?|  	�5 A|  *�N  F	�Ze     +*	 I@   	�Ze     *0O  M	��e     *<O  N	�Ze     +�Z Q@   	Ef     +�Y T@   	Ef     +*\ W@   	xDf     +�X Y	�   	PEf     +q\ \@   	hDf     +w\ ]@   	pDf     +�\ ^@   	�Df     +�V a|  	tDf     +"W crH  	`Df     �   �P  9   9    +�V e�P  	 Ze     +xX o@   	HEf     +�Z p@   	�Df     + Y q@   	Ef     �   Q  9    +�[ s�P  	0Ef     + u|  	|Df     */M  v	Ef     	P! {|  �   lQ  9   	9    +$Z |VQ  	`Ef     �   �Q  9   � +_[ ~�Q  	`Ff      �	�Q  �f  �E   � �
�Q  KZ �rH  �\ �
�    �   �Q  9   	 �[ ��Q  i[ (�gR  �\ �E   gW �gR  �\ �mR  KZ ��	  x �E   y �E  "\ �E  $ R  �Q  p[ �R  +�W �E  	�Df     +:W �E  	(Ef     +8Y �E  	�Df     �   �R  9    +�Y �
�R  	 Ze     +jV �	�R  	 Ef     sR  
W   �<S    ޽  :	  Y 1W [  +�Z �S  	�Df     �Q  bS  9    +G] �RS  	@Ye     +�\ �	sR  	 Ye     #W   �S  ,ep1  ,ep2 ,ep3 ,ep4 �Y  -Y �S  	�Df     �Q  �S  9    -=[ �S  	�Xe     -�V 	sR  	@Xe     #W   *ET  W  pW W �W ��  JV  -3[ 1T  	 Gf     �Q  lT  9    -CY 3\T  	�We     -:] <	sR  	`We     #W   L�T  �p   +�  ��  �Z �X �V �W �\ [  -4Z V�T  	Ef     �Q  U  9    -.X X�T  	`Ve     -�\ d	sR  	 Ve     #W   rQU  [  �V  -�Z u5U  	 Ef     �Q  xU  9     -�Y whU  	 Ve     -ZY |	sR  	�Ue     #W   ��U  �V  lY  -hX ��U  	XEf     -�Y �hU  	�Ue     -cY �	sR  	`Ue     #W   �5V  �W  \W �X vY Y  -pX �V  	Ef     -.Y ��S  	�Te     -Z �	sR  	�Te     #W   ��V  _\  �\ �\ e\ �\ k\ Z  -GX �zV  	�Df     -�Y �RS  	�Se     -'] �	sR  	�Se     -�V �RS  	�Re     -] �	sR  	�Re     �   7W  9   O -�X �	'W  	�Df     .epi �	@   	lDf     /X ��R  	�B     /�X ��R  	ЧB     -vV Q		  	�Re     -�W ]		  	`Re     0� �@     �       �0�  ۲@     '       �1�[ ��@            �&X  2W[ �R  U 3uZ �4�  ���@     �      ��Y  5x �E  	��e     5y �E  	��e     6i �W   �  �  6max �W   ��  ��  /b[ �'W  ��7� ��   ��  ��  7' �@   ��  ��  8@  cY  7>Z �
@   o�  k�  9��@     y  Y  :Uw :QP 9��@     y  6Y  :Uw :QP 9Ц@     3`  NY  :Uw  ;��@     �^  :Qw   <,�@     �_  9z�@     y  �Y  :T8 <��@     y  9��@     y  �Y  :T8 <�@     y   3�  k= e  �	|  �@     	      ��^  >ev ��^  ��  ��  6ch �@   	�  ��  6key �@   D�  .�  6i �@   6�  0�  /�Z �@   	 �e     /�Z �@   	��e     /�" �@   	��e     /?\ �@   	��e     /�" �@   	��e     /9\ �@   	��e     ?&X  �@      �@     
       6@�^  c�@       c�@            L[  A�^  ��  �   <!�@     &y  <U�@     +e  9r�@     2y  N[  :U0:TG 9y�@     Ud  e[  :U0 <��@     >y  <��@     >y  <ک@     >y  <��@     >y  <�@     >y  <@�@     >y  <]�@     >y  <��@     >y  <��@     >y  <��@     >y  <$�@     >y  <S�@     >y  <o�@     >y  9�@     y  2\  :T	0Ef     :QH <A�@     �l  <U�@     Jy  9��@     3`  d\  :Us  B�@     x\  :Us  <2�@     Vy  <��@     �c  <��@     �Y  <í@     �Y  9ϭ@     2y  �\  :U0:TG 9֭@      l  �\  :U0 <�@     �Y  9��@     2y  ]  :U0:TG 9��@     Hm  ]  :U0 <�@     �Y  95�@     �c  C]  :U0 9N�@     2y  _]  :U0:TG <S�@     �k  9l�@     2y  �]  :U0:TG 9s�@     f  �]  :U0 9��@     Wf  �]  :Uu  9��@     2y  �]  :U0:TG <��@     �k  9��@     y  ^  :U	�RB     :T8 <�@     by  <�@     �Y  9Y�@     2y  :^  :U0:TC 9��@     2y  V^  :U0:TC 9�@     2y  r^  :U0:TF 9m�@     2y  �^  :U0:TF Bܰ@     �^  :U1 ;ѱ@     2y  :U0  �  C�W {|  �^  Dkey {@    1�[ MH�@     n       ��_  >x N@   ��  ��  >y O@   ��  ��  Eb[ P
�   7�  3�  6w R
@   v�  p�  6ch S�   ��  ��  6c T
@   �  �  6cx U
@   h�  \�  6cy V
@   ��  ��  <}�@     Jy  ;��@     y  :U~ :Tv   FZ :@   �@     :       �3`  Eb[ :�   &�  $�  6i <-   M�  I�  6h =@   ��  ��  7  >@   ��  ��   FNX #@   ��@     Q       ��`  Eb[ #�   ��  ��  6i %-       6w &@   �  �  6c '@   �  �  <�@     Jy   0�Z ��@            �1$[ 	A�@     5       �a  2b[ 

�   U2KZ 
G   T2�X |  Q 1SV ��@     4       ��a  E��   �R  �  �  E�[ @   N H 9'�@     y  �a  :U	��B     :T8 GA�@     y   1�\ �١@     4       �b  E��  ��R  � � E�[ �@   � � 9�@     y  b  :U	��B     :T8 G�@     y   1:X ��@     �       ��c  >x �@   H > >y �@   � � E�Y �@   ) # E�X �@   { u 6xx �
@   � � 6i �
@   � � 9�@     y  �b  :U	m�B     :T8 9#�@     y  �b  :Usx:T|  9:�@     y  c  :U	v�B     :T8 9L�@     y  *c  :Ux:T|  9g�@     y  Nc  :U	�B     :T8 9w�@     y  lc  :Uv :T|  9��@     y  �c  :U	��B     :T8 H��@     y  :U�R3$�U"#:T�T  1] �,�@     R       ��c  E�W �@   � � G~�@     ny   1�W �ל@     U       �9d  E�W �@   ' # <��@     ny   I�Y �Ud  J�W �@    1T\ ��@     Y       �e  E�W �@   b ^ Ke  �@      �  ��d  L�  Me  � �   9X�@     zy  �d  :U	`Ff     :T�:Q	��B      Hm�@     �`  :Uu :Tt :Qq   C�Z {�   +e  N_�  }1B   I�W kGe  Dkey k@    IKW Ece  J�W E@    1�[ 3��@     !       ��e  E�W 3@   � � OGe  Ѳ@      Ѳ@     
       A	AUe  � � G۲@     �W    1/] -��@     
       �f  E�W -@   ' # H��@     �W  :Uu   I�W ;f  J�W @    I\ Wf  Dkey @    1X ��@     K       ��f  E�W �@   b ^  1�Y ���@     
       ��f  E�W �@   � � H��@     �W  :Uu   1�[ ��@     �       ��g  9�@     y  g  :U	��B     :T8 9(�@     y  5g  :Ul:T? 9A�@     y  Lg  :T8 <`�@     y  9y�@     y  pg  :T8 <��@     y  9��@     b  �g  :Q: H١@     b  :Q9  I\ ��g  J�W �@    IgZ ��g  J�W �@    I�Z ��g  Dkey �@    1�V �ߚ@     #       �Zh  9�@     y  ?h  :U	�B     :T8 H�@     y  :U6:T&  I�Y �vh  J�W �@    1�[ ���@     D       �i  9��@     y  �h  :U	��B     :T8 9��@     y  �h  :U`:T> 9̚@     y  �h  :U	�B     :T8 Hߚ@     y  :U6:T&  1A] zx�@     #       �ri  9��@     y  Xi  :U	��B     :T8 H��@     y  :U^:T2  1�Y c��@     7       ��i  E�W c@   � � Gל@     �y   1�[ Ri�@     7       ��i  E�W R@     G��@     �y   1�Y M �@     
       �?j  E�W M@   N J H
�@     �W  :Uu   1�V B��@     f       ��j  9��@     y  �j  :U	��B     :T8 9 @     y  �j  :U<:T& 9�@     b  �j  :Q@ H�@     b  :Q@  1�X 4Q�@     '       �'k  9k�@     y  k  :U	�B     :T8 Hx�@     y  :U0:T0  1�X ���@     �       ��k  7� ��   � � 7w[ �	@   � � 7~[ �@     9�@     �y  �k  :U	$�B      9K�@     y  �k  :T8 ;W�@     y  :U0:T0  3\X �IyW ��k  Dkey �@    3�\ �ISZ � l  Dkey �@    IW �<l  J�W �@    1�V {8�@     i       ��l  E�W {@   I C 9k�@     y  �l  :U	0Ef     :Tv :QH ;x�@     �y  :Uv :T	�B       1aV n��@     4       �.m  E� n@   � � P&X  ��@      @  q;��@     �y  :Us :Ts H`Ef     "  IOY YHm  Qi [@    IX Idm  J�W I@    1}\ <�@     6       �n  E�W <@   � � /� >n  ��}?&X  &�@      &�@     
       C9�@     �y  �m  :U�U 9�@     y  n  :Uw :Q
  ;&�@     �y  :Uw   �   )n  9   � 1�Z %"�@     p       �9o  >x %@   8	 ,	 >y %%@   �	 �	 Qi '@   9C�@     y  �n  :U	R�B     :T8 9P�@     y  �n  :Usx:Tv  9_�@     y  �n  :U	[�B     :T8 9n�@     y  �n  :Usx:Tv  9��@     y  !o  :U	d�B     :T8 H��@     y  :T�T#  1] ��@     h       ��o  Qi @   9Ϥ@     y  �o  :U	�B     :T8 9�@     y  �o  :UH:TL <��@     )n  ;�@     �^  :Qvh  1�V �v�@     �       ��p  7t �  D
 <
 6i �@   �
 �
 /� �n  ��}9��@     �y  6p  :Us  9��@     y  Up  :Uw :Q
  9��@     �y  zp  :Uw :T	P�B      9ƞ@     y  �p  :Uv :T	�B     :QH 9�@     �y  �p  :Uv :T1:QH:R|  ;��@     �y  :U|   R9d  ~�@     +       �-q  AGd  �
 �
 S9d  ��@            AGd  . ,   R+e  ��@     S       ��q  A9e  Z R T+e  `  A9e  � � 9�@     2y  �q  :U0 9�@     �y  �q  :Ui G��@     &y    R�k  ��@     "       �r  A�k    T�k  �  A�k  g c <�@     dm  H�@     2y  :U0:TH   R�g  �@     .       ��r  A�g  � � T�g  �  A�g  � � ?&X  ?�@      ?�@     
       �;?�@     
z  :U4:Q1   R;f  L�@     *       ��r  AIf  5 / S;f  T�@     !       AIf  � � P&X  p�@        Gu�@     z    Rl  Ɵ@     "       �^s  Al  � � Tl  p  Al    <ڟ@     �l  H�@     2y  :U0:TH   R�k  v�@     a       ��s  9¢@     zy  �s  :U	�Df     :TP:Q	�B      Gע@     �`   Rf  ע@     =       �/t  A-f  Q M Uf  �@            !t  A-f  � � H�@     2y  :U0:T"  G�@     �`   R�g  m�@     9       ��t  A�g  � � U�g  r�@            �t  A�g  1 / H��@     �`  :Uu :Tt :Qq   ?&X  ��@      ��@     
       �;��@     
z  :Q1  R.m  �@     �       ��u  V<m  8   4u  M<m  W U <��@     3`  Hǥ@     �^  :Q	-�B       97�@     y  Xu  :U	%�B     :T8 9I�@     y  uu  :UH:TL <^�@     )n  ;}�@     �^  :Qvh  W�Y  ˥@     ,       �W&X  �@            �RHm  �@     (       �Zv  AVm  � z UHm  �@            4v  AVm  � � H#�@     �`  :Uu :Tq :Qq   9.�@     �W  Lv  :Uu  G4�@     �o   R l  4�@     2       ��v  A.l  + ! U l  =�@            �v  A.l  � � HK�@     �`  :Uu :Tq :Qq   9_�@     �W  �v  :Uu  Ge�@     �o   R�k  f�@     �       ��w  X{�@     2y  'w  :U0:T" <��@     �Y  <��@     �o  9��@     �W  Yw  :Uu  9Ѩ@     zy  �w  :U	�Df     :TP:Q	��B      H�@     �`  :Uu :Tt :Qq   RZh  
�@     A       �)x  Ahh  � � UZh  �@            x  Ahh  K G H*�@     �`  :Uu :Tq :Qq   GK�@     �W   R�g  K�@     Q       ��x  A�g  � � U�g  Z�@            �x  A�g    ;h�@     �`  :Uu :Tq :Qq   9��@     "z  �x  :U	k�B      G��@     �W   RGe  ��@     
       �y  AUe  E A H��@     �W  :Uu   Y  /'	Y��  ��  CY� � ?Y/ / 05Y� � +6Y  1Y� � 2Y�/ �/ %HY� � hY�[ �[ �Y[�  [�  fY�X �X +SYE\ E\ +TY��  ��  07Y'�  '�  3Y�$ �$ %1Y� � (#Y� � %,Y�/ �/ [Y�K �K �Y5L 5L YYsK sK 1'Y� � %&Y� � 
(Z�E �E 4  �   �P  S#  �^ �*  ��@     �      � �d  �)  �=   ,	  ^&  nC (W   �E `   p   p   =     D  �   �E  �    �G  �   F  �   3E  �    �  	
�1  @9  Q  9   �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2K  8;:  5K  < ?  1  ?  int �K 8"�   �  Kj  R  �  Lj  �  Mj  9�  uO 	K  YP 9  kS 9  e2  0t  �    �0  }  ��  �  �   	J  D   �C  
D  ���� �C  	N�  ڵ  	R�    ��  
�9  �\  
�  �  
�M  �  ��  
�K  ��  
�K  2�  
�  ��  
�K  Ɇ  
�#  ��  
�K  ��  
�K  �h  
�K  rK  
�K  l�  
�K  ]�  
�K  ��  
�K  *  cK   K     =    N�  %�  ��  '#  =� $  
��  .Y  ^�  2�   }�  7#  �� ;�    	�  r�  �   .� $�  O� )�   �  �  9     �  �  �   �  1   �  �  �   �   1    �  ��  ,Y  �  oS  '�  
dS  ()T  � +
T   � ,�  @�  -
K  >z .
K  �  /�   �H  3d    ?  d  =    �  �� 7d  �� 8�   �   "�  ��  WH  �~  �O  �m  ��   �  ��  ��  	 G�  �K  �@     �       �d  buf �9  � | �a �"1   � � s �7d  � � �L ��  ��~��  �	K  5 3 ��@     j  R��~  F  �F �K  �   buf �9  !�a �#1    s �8d  !�L �C�  "��  �	K   p   ��  �9  ��@     $      ��  s � d  Z X ��  �9  � } #v �d  �L ��  ����  �1   � � $I�@       W  Us  $]�@       v  U	��B      $m�@       �  Uv T| Qs  ù@     ~  Uv Qs   �	 �	  k�@     B       �  s �&d    ` �5d  B @ ��@     %  T�T  �` �	  *�@     A       �~  s �(d  g e ? �7d  � � ^�@     1  U�UT�T  ` �	  �@     $       �  `5 �9  � � src �0d  � � �_ �<1     82  �1   R N %*�@       T�T   u	  R  !`5 u9   src u.d  !�_ u:1   #len w1    t] 79  �@           ��	  �a 7#d  � � &_ 79d  � � P] 8#d    ��  :9  N H &dst :9  � � &p ;d  � � �_ <1   L J ��  =1   q o 
^ =1   � � $Q�@     =  H	  T~  $|�@       `	  Us  $��@       	  U	m�B      $��@     1  �	  Uv T~ Q|  ��@       U Tw Qs   aa $9  ��@     9       �F
  ` $%d  � � ��  &9  %  $��@     I  *
  Us  ��@       U	E�B       �` 9  �@     t       �  �a 9  p n &_ *9  � � �^ �   � � �_ �   � � &len �     &i �   @ < p�@     U  U| T~ Qs   '�` ���@            �X  (� �9  { w )p �9  � � *�@     a   '�^ ���@     u       �
  (�> �9    (`5 �*9  6 * )src �9  � � +��  �9  o g +�� �	K  � � *ȵ@     a  %��@     m  U	�B     Q�T  ,SJ �	  �@     m       ��  -str � d  M G (��  �*�  � � $5�@     y    Us T	�B     Qv  $R�@     y  �  Us T	�B     Qv  $h�@     y  �  Us T	�B     Qv  ~�@     y  Us T	��B     Qv   K  ,>1 �9  ѹ@            ��  -s �9     .f` �9  
ɨB     �%�@     �  U	ɨB     T	(�B     Q�UR0  ,�_ �K  ��@     �       �  (� �9  X R (�< �#  � � +t �j  � � +r� �	K  2 0 +�� �K  W U )buf �#  � z $��@     �  B  U| T	P�B      $��@       g  U	�B     T|  $ƴ@     �    Uv  $״@     �  �  T1Q0 $�@     �  �  U} T1Qs  $ &Rv  $��@     �  �  Uv  �@       U	�B     T|   #  ,�. p	  D�@     H       ��  (� p9  � � (m�  p'�   $  (�� p3K  v p +t rj  � � +r� s	K  � � $W�@     �  �  U�UT	��B      $t�@     �  �  U| T1Qv  $ &Rs  �@     �  Us   ,�] ZD   �@     >       ��  (t Zj  '  !  +�_ \
D   w  s  +�� ]
D   �  �  $�@     �  p  Us  $$�@     �  �  Us T0Q2 $,�@     �  �  Us  <�@     �  Us T| Q0  ,$�  B	  ȳ@     >       �H  (��  B9   ! �  +}_ Dj  =! 9! $ӳ@     �  :  U�UT	w�B      *�@     �   'xT 7��@     
       ��  (�> 79  w! s! %ȳ@     �  U�UT
�  /  Ƕ@     >       �?  0  �! �! 0*  
" " 07  q" i" 1D  2  �  37  0*  �" �" 0  &# "# 4�  5D  c# _# �@     �  U�UTs Q�Q1    /j  �@     /       �  0|  �# �# 0�  $ $ 0�  t$ n$ 0�  �$ �$ 1�  2j  �  0�  % % 0�  S% O% 0�  �% �% 0|  �% �% 4�  5�  2& 0& ��@     �  Uv Ts Q�QR�R    6��  ��  A6��  ��  76'�  '�  6-` -` 6�` �` (6��  ��  	6� � 6� � 6��  ��  d6�Q �Q h6�/ �/ [6� � 66�K �K �65L 5L Y6�L �L �6pL pL �6VL VL �6�^ �^ 6�` �` 6�F �F m �    �S  S#  b �*  ��@     G       � Jh  T   A   F   � 1   ,	  e2  M    b A   	�B     *b .�   	�e     int )b /�   	�e     	�( >Һ@            �
� 8�   ��@            �
� 2�   ��@            � �O   <T  S#  �b �*  �@     B      x [h  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  
K   "f  ��  WH  �~  �O  �m  ��   �  ��  ��  	 0t  r  e2    �0  }  ��  f  
K   J�  D   �C  
D  ���� �C  N�  ڵ  R�  �  
K   &  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
K   /_  ��   [r  �4 #�  �   �X  52  
K   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  Kk  
�   P  =_  ��   R�  N�  ��  ��   �p  W�  
K   	3@  ��   ({  ��  ğ   F]  	8  
K   	Y�  ��   �c  |  ��  l  ��  �   
K   	k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  	{�  
K   	�  &�   �  º  GY  �f  ��   v�  	��  
K   	�Z  GQ   ϼ  �  �_  X  &�  �b   t�  
 �   Z  f  |  =   �' k  	��  1|  	]  4�  f  f  �  =   � �  	Zy  8�  �  �  =   =   � �  	��  ;�  Ʃ  QK   �  �  
  =     �  	�  W
  �p  #'  -  4   S�  $@  F  Q  R    T}  %]  c  s  R   R    '	�  acv )  ��  *4  ��  +Q   �y -s  �Y  6�  ��  :�  s�  <�   �H  =�  xz  >�   �  x @�  �    =    y     =    
�	g  x ��   y ��  Mp ��  *� ��  ޽  ��   ~x �   
K   �	  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �s  
K   �W#  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�	  (x	�#  �u z�	   � {	�   s |	�   � ~�  N�  W#  ��  �	�   ��  �	�     J]  �d#  �#  �#  =   � �^  ��#  �   $    �  ��#  !K   �`'  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  $  \	�(  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /m'  �(  �(  =   � ��  1�(  �]  ���*  `e ��   x �Z  y �Z  z �Z   ��  ��*  (cN  ��*  0Mp ��  8�u ��	  <� ��   @�H  ��*  Hr�  ��*  P��  ��*  X��  �Z  `m�  �Z  d��  �Z  h  �Z  l3F  �Z  p8F  �Z  t=F  �Z  x��  ��   |*� �`'  �y� ��*  �s ��   ��� �+  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  �*  ���  �   ���  	�   ��R  �,  �f�  �   �I}  g  ���  �*  � �(  Gx  ��*  >} �E0   �}  ��  �|  ��  
 �*  �(  �#  "d  HN�,  mo P�.   ��  Q�6  cmd Re6  �  WZ  (_  YZ   #_  [Z  $bob ]Z  (�  a�   ,�[  b�   0sb  d�   4d]  g�6  8�W  h�6  P��  i�  h�� l/  l�N  m�  |E�  p�  ��W  r�6  �~�  s/  �*� t/  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��.  �#�R  ��    #��  ��   #�  ��   #h  ��6  #I�  ��  @ +  �z �(  �  	��  ��   	�\  ��  	�  �-  �  	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  ��,  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	�-  x EZ   y FZ   �{ H�-  (T	.  `e V�   x WZ  y XZ  z YZ    	�  [�-  �a	�.  = cZ   F�  dZ  �~ e�  h�  f�  
t�  g�  �k h�  tag i�  �N  l
�   ��  o�.  ��  r
/   iK  u.  0��  x
�   XS�  {�.  `��  ~R   h��  ��   pu| ��/  x �,  �   /  =    �}  X��/  v1 ��0   v2 ��0  dx �Z  dy �Z  �  ��  �k ��  tag ��  �W  �   �o ��0  $��  �~0  4SX  �E0  8d�  �E0  @��  �
�   H��  �R   P �/  /  �z �%.  �	E0  2�  �Z   ]  �Z  �h  ��  �N  ��  
�K  ��  >} �E0   �/  �}  ��/  
K   �~0  ��   �  o�  ��   ��  �W0  �-  Z  �0  =    �u  �/  �z ��*  8�	(1  v1 ��0   v2 ��0  82  �Z  Mp ��  [�  �(1   �  �.1   SX  �E0  (d�  �E0  0 K0  �0  A{ ��0  4	�1  $x Z   $y 	Z  $dx 
Z  $dy Z  �o �1  )�    0 Z  �1  =   =    (} @1  �  *�  %v  @2~2  @�  4~2   $x1 5�   $x2 6�   .]  8Z  5]  9Z  �� :Z  ��  =�   �  @Z   ��  CZ  $�n  G�2  (9x  H�2  0�^  I�2  8 41  �  >�  K�1  %�h  PRs3  s�  Us3   �H  Vs3  $x1 X�   $x2 Y�   $gx \Z  $gy ]Z  $gz `Z   $gzt aZ  $�x  dZ  (� fZ  ,~�  iZ  0t  kZ  4.� l�   8�  py3  @	�  r�   H �2  �1  �h  t�2  �	�3  �c  ��   �O  ��3  �x  �
�3   �  �3  =    �  �3  =    I�  ��3  �	4  �  ��    �  �4   �3  �  ��3  &��	�4    �Z   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  $top �	�4  '��  �	�  U'��  �	�  V'� �	�4  W'�  �	�  � �  �4  =   ? ��  �(4  	H5  ~�     �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�4  H5  d5  =    	S�  'T5  
K   7�5  {�   U�  ~�   >	�5  �� @+   s A
�   sx BZ  sy CZ   Nz E�5   	e6  ��  "�   E�  #�  e% $�  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�5  
K   1�6  ��   ��  ��   �y  9q6  �   �6  =    �  �6  =    �  �6  =    �5  �6  =    hy �+  (�	N7  in ��   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
/  �a  �
�   $ ��  ��6  ��	�7  2�  �
�    I�  ��  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��7  ( N7  8  =    ޴  �Z7  	.L  &8  Z  	׮  )8  	�  +8  	�  ,8  	�Q  .y3  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�8  �   	��  8�8  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�8  4  	��  H�   	��  I�0  	��  K�   	a� L~2  	w�  N�   	P{ OE0  	��  Q�   	��  RA9  �0  	��  T�   	�� U_9  �1  	�}  W�   	u| X.1  	M�  Z�   	P�  [(1  	��  aZ  	��  bZ  	�  cZ  	�p  e�  	�T  f�9  �6  	�a  j�  �   �9  =   � 	ը  l�9  �  :  =   @ 	�p  m :  	 �  pZ  	p|  q�  	$Y  v�   	�K  y�   	g  {Y:  �4  	d�  |Y:  	��   Z  		�  !Z  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +Z  	`�  ,Z  	A�  -Z  	��  /�   	��  1�   	P�  2�   y3  ;  =   =   / 	��  E�:  y3  -;  =   / 	Ԁ  F;  y3  O;  =   =    	7� G9;  	�R  I�   	��  Jy3  	��  U�   (	P�  \�;  ;  	��  ]�;  	L�  ^�;  	ߵ  _�;  	�  a�;  	@�  ~2  	[�  (1  	 �  .1  	SX  E0  	d�  E0  	��  �   	_�   �   	��  "�  	��  %�  	'�  &�  	�]  (�  �2  V<  =   � 	�P  *F<  	ӯ  +n<  �2  	|  -�<  y3  	��  .�<  	��  /�<  �<  �<  �   �    	��  �2  �   �<  	qY  "�<  	�  #�<  �  �<  =   ? 	��  %�<  	��  &�<  Z  =  =   � 	@Y  (=  Z  :=  =   ? 	V�  ))=  3  V=  =    	�h  F=  	�  n=  3  	�  3  	�f  !�<  	r�  "�<  	��  %�2  	��  &�2  	׆  'Z  	��  (Z  	�  *Z  	��  +Z  	�  y3  	��  �   	�_  �   	�_  �   	b  Z  	t  Z  	j�  "�,  	�  :�   	��  ;�   	��  <�   	�W  >y3  	hn  @Z  	U~  AZ  	�  BZ  	 �  CZ  	%�  F�,  	�u  H�,  	z  I�,  	ʓ  C�  g  �>  =    	��  b�>  �   �>  =    	��  c�>  	0K  d�   	?�  e�   �	L?  x �Z   y �Z  dx �Z  dy �Z   ��  �?  �z?  �p �
�.  ��  �
.1   �	�?  {q �Z   ��  ��  d �	X?   t�  �z?  �?  �?  =   � 	r ��?  	�T  ��?  �?  	l�  �Z  	�  �Z  	?k  �Z  	�d  �Z  	2~ �L?  	��  ��  	��  �Z  	k�  �Z  	Z�  �.1  .1  _@  =    	�v  �O@  	�v  ��   	"�  ��.  �  �,  �U  �2  ��  �2  t�  �   �  	�   .Y  
Z  7Y  Z  �h  �@  �.  *� /  <i  /  	G  �  	��  �   �   3A  =    
K   �TA  )top  �G  �  �]  �3A   �	�A  ��  �.1   ��  �TA  O{  �
�   ��  �
�   iK  ��A   .  ��  �`A  �A  �A  =    	��  ��A  !K    B  )up  �  �F  �S   FT  
�A  !K   ;B  ��   �x  H�  ��  �H   ��  B  H	�B  `e �   >} E0  L� Z   $low Z  $+�  Z  (�Z !
�   ,r� "
�   0�f  # B  4�f  $ B  8��  %�  <$tag &
�   @*� ';B  D �w )HB  C  C  =    �B  �  2C  !K   �_C  ��   �s  z�  ��  �T  ܭ   gY  �+C  H�	D  `e ��   *� �_C  >} �E0   �W  �Z  (�}  �Z  ,L� �Z  0��  ��  4��  �
�   8$tag �
�   <��  �
�   @  w �lC   D   D  =    D  j�  D  !K   XTD  )ok  �b �b  Mb ]3D  ) mD  J @�D  � "�    � '
#A  �� *	�   
 -�D  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 aD   H	AE  � K�    C� N	�   "8 QR   t TR    . VE  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   aD  �E    	R �E  AE  �E    	� �E  
K   rfH  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	  V�   e6  	��  !M�  	(h  !N�   	l�  !N�   	�  ".�  	�  "/�  	�  "0�  	�  "2�  	w�  "8_  	�  "9&  	�  ":�  	�_  ";�   	��  ">�  	�  "J�  	"�  "R  	t�  "S�   	�w  "T�   	؜  "Y�   	q�  "[�  	Ƚ  "^  	�  "_�   	�y  "`�   	b�  "c�   	+�  "f�  	��  "i�  	֘ "l�   	�J  "x�   	��  "y�   	ks  "�   	�  "��   	J�  "��   	�i  "��   	��  "��  	��  "��  	��  "��  	<� "��  	��  "��  	��  "��  	5�  "��  	<m  "��   	 K  "��   	�R  "��   	op  "��   	�m  "��   	D  "��   	X�  "��   	If  "��   	� "��   	��  "��  	�U  "��  	`  "��  	J�  "��  	��  "��  	� "�@  �6  K  =    	�  "��J  �   K  =    	� "�K  g  <K  =   	 	,�  "�,K  	R�  "�TK  g  g  jK  =    	�u  "�ZK  	��  "�8  	�e  "��   �   �K  =   � 	(�  "��K  	�  "��  ��  "@  �v  "�   n�  "�   4�  "�   *b "�   ��  "rH  *&D  &	 Gf     +�b /�   �@     B       �rL  ,��  /!.1  U-i 1
�   [& U& -rtn 2
�   �& �&  .�b ��@     6       ��L  ,��  (.1  U-i 
�   �& �&  .�b 	�@     :       �M  /c ' D  Q' I' -i 
�   �' �' 0*�@     nO  1U�U  2�b ��@     "       �LM  3c �$ D  U4i �
�   7( 1(  5@b ��   ��@     &      ��N  6��  �.1  �( �( 6*� �_C  �( �( 7�k �
�   3) ') 4rtn �
�   �) �) 4sec �E0  4* 2* 7�x � D  ]* W* 8߼@     rL  �M  1Uu  8��@     zO  N  1U~ 1T}  8+�@     �O  >N  1UH1T61Q0 86�@     �O  VN  1Us  8��@     �O  nN  1Uv  0Խ@     M  1Uu   2c -C�@     H      �nO  6�x -  D  �* �* 4res /TD  J+ :+ 8x�@     �O  �N  1R01X1 8��@     �O  �N  1TF 9ʻ@     �L  O  1U�U 8�@     �O  ,O  1TC 8	�@     �O  CO  1X1 8,�@     �O  ZO  1TF 0X�@     �O  1TC  :c c H:Vb Vb `:� � 6:3b 3b G:nb nb ]	;c c `:� �  6 nR   �W  S#  ?c �*  )�@     �      ! �j  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  
K   "f  ��  WH  �~  �O  �m  ��   �  ��  ��  	 0t  r  e2    �0  }  ��  f  
K   J�  D   �C  
D  ���� �C  N�  ڵ  R�  �  
K   &  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
K   /_  ��   [r  �4 #�  �   �X  52  
K   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  Kk  
�   P  =_  ��   R�  N�  ��  ��   �p  W�  
K   	3@  ��   ({  ��  ğ   F]  	8  
K   	Y�  ��   �c  |  ��  l  ��  �   
K   	k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  	{�  
K   	�  &�   �  º  GY  �f  ��   v�  	��  	"|  
*�  	��  
+�  	I�  
,�  	�a  
-�  t�   �   Q  ]  s  =   �' b  	��  1s  	]  4�  ]  ]  �  =   � �  	Zy  8�  �  �  =   =   � �  	��  ;�  Ʃ  QK   �  �    =     �  	�  W  �p  #  $  +   S�  $7  =  H  R    T}  %T  Z  j  R   R    '	�  acv )  ��  *+  ��  +H   �y -j  �Y  6�  ��  :�  s�  <�   �H  =�  xz  >�   �  x @�  �    =    y    =    
�	^  x ��   y ��  Mp ��  *� ��  ޽  ��   ~x �  
K   �	  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �j  
K   �N#  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�	  (x	�#  �u z�	   � {	�   s |	�   � ~�  N�  N#  ��  �	�   ��  �	�     J]  �[#  �#  �#  =   � �^  ��#  �   �#    �  ��#  !K   �W'  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  $  \	�(  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /d'  �(  �(  =   � ��  1�(  �]  ���*  `e ��   x �Q  y �Q  z �Q   ��  ��*  (cN  ��*  0Mp ��  8�u ��	  <� ��   @�H  ��*  Hr�  ��*  P��  ��*  X��  �Q  `m�  �Q  d��  �Q  h  �Q  l3F  �Q  p8F  �Q  t=F  �Q  x��  ��   |*� �W'  �y� ��*  �s ��   ��� ��*  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  �*  ���  �   ���  	�   ��R  �,  �f�  �   �I}  ^  ���  �*  � �(  Gx  ��*  >} �<0   �}  ��  �|  ��  
 �*  �(  �#  "d  HN�,  mo P�.   ��  Qh6  cmd R;6  �  WQ  (_  YQ   #_  [Q  $bob ]Q  (�  a�   ,�[  b�   0sb  d�   4d]  gt6  8�W  h�6  P��  i�  h�� l�.  l�N  m�  |E�  p�  ��W  r�6  �~�  s�.  �*� t�.  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��.  �#�R  ��    #��  ��   #�  ��   #h  ��6  #I�  ��  @ �*  �z �(  �  	��  ��   	�\  ��  	�  �-  �  	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  ��,  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	�-  x EQ   y FQ   �{ H�-  (T	.  `e V�   x WQ  y XQ  z YQ    	�  [�-  �a	�.  = cQ   F�  dQ  �~ e�  h�  f�  
t�  g�  �k h�  tag i�  �N  l
�   ��  o�.  ��  r
�.   iK  u.  0��  x
�   XS�  {�.  `��  ~R   h��  ��   pu| ��/  x �,  �   /  =    �}  X��/  v1 ��0   v2 ��0  dx �Q  dy �Q  �  ��  �k ��  tag ��  �W  ��  �o ��0  $��  �u0  4SX  �<0  8d�  �<0  @��  �
�   H��  �R   P �/  /  �z �.  �	<0  2�  �Q   ]  �Q  �h  ��  �N  ��  
�K  ��  >} �<0   �/  �}  ��/  
K   �u0  ��   �  o�  ��   ��  �N0  �-  Q  �0  =    �u  �/  �z ��*  8�	1  v1 ��0   v2 ��0  82  �Q  Mp ��  [�  �1   �  �%1   SX  �<0  (d�  �<0  0 B0  �0  A{ ��0  4	�1  $x Q   $y 	Q  $dx 
Q  $dy Q  �o �1  )�    0 Q  �1  =   =    (} 71  �  *�  %v  @2u2  @�  4u2   $x1 5�   $x2 6�   .]  8Q  5]  9Q  �� :Q  ��  =�   �  @Q   ��  CQ  $�n  G{2  (9x  H{2  0�^  I{2  8 +1  �  >�  K�1  %�h  PRj3  s�  Uj3   �H  Vj3  $x1 X�   $x2 Y�   $gx \Q  $gy ]Q  $gz `Q   $gzt aQ  $�x  dQ  (� fQ  ,~�  iQ  0t  kQ  4.� l�   8�  pp3  @	�  r�   H �2  �1  �h  t�2  �	�3  �c  ��   �O  ��3  �x  �
�3   �  �3  =    �  �3  =    I�  ��3  �	4  �  ��    �  �4   �3  �  ��3  &��	�4    �Q   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  $top �	�4  '��  �	�  U'��  �	�  V'� �	�4  W'�  �	�  � �  �4  =   ? ��  �4  	?5  ~�     �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�4  ?5  [5  =    	S�  'K5  >	�5  �� @�*   s A
�   sx BQ  sy CQ   Nz Eg5   	;6  ��  "�   E�  #�  e% $�  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�5  
K   1h6  ��   ��  ��   �y  9G6  �   �6  =    �  �6  =    �  �6  =    �5  �6  =    hy ��*  (�	$7  in ��   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�.  �a  �
�   $ ��  ��6  ��	�7  2�  �
�    I�  ��  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��7  ( $7  �7  =    ޴  �07  	.L  &�7  Q  	׮  )�7  	�  +�7  	�  ,�7  	�Q  .p3  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7c8  �   	��  8c8  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�8  4  	��  H�   	��  I�0  	��  K�   	a� Lu2  	w�  N�   	P{ O<0  	��  Q�   	��  R9  �0  	��  T�   	�� U59  �1  	�}  W�   	u| X%1  	M�  Z�   	P�  [1  	��  aQ  	��  bQ  	�  cQ  	�p  e�  	�T  f�9  �6  	�a  j�  �   �9  =   � 	ը  l�9  �  �9  =   @ 	�p  m�9  	 �  pQ  	p|  q�  	$Y  v�   	�K  y�   	g  {/:  �4  	d�  |/:  	��   Q  		�  !Q  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +Q  	`�  ,Q  	A�  -Q  	��  /�   	��  1�   	P�  2�   p3  �:  =   =   / 	��  E�:  p3  ;  =   / 	Ԁ  F�:  p3  %;  =   =    	7� G;  	�R  I�   	��  Jp3  	��  U�   (	P�  \b;  U;  	��  ]b;  	L�  ^b;  	ߵ  _b;  	�  ab;  	@�  u2  	[�  1  	 �  %1  	SX  <0  	d�  <0  	��  �   	_�   �   	��  "�  	��  %�  	'�  &�  	�]  (�  �2  ,<  =   � 	�P  *<  	ӯ  +D<  �2  	|  -V<  p3  	��  .V<  	��  /V<  z<  �<  �   �    	��  {2  �   t<  	qY  "�<  	�  #�<  �  �<  =   ? 	��  %�<  	��  &�<  Q  �<  =   � 	@Y  (�<  Q  =  =   ? 	V�  )�<  v3  ,=  =    	�h  =  	�  D=  v3  	�  v3  	�f  !�<  	r�  "�<  	��  %{2  	��  &{2  	׆  'Q  	��  (Q  	�  *Q  	��  +Q  	�  p3  	��  �   	�_  �   	�_  �   	b  Q  	t  Q  	j�  "�,  	�  :�   	��  ;�   	��  <�   	�W  >p3  	hn  @Q  	U~  AQ  	�  BQ  	 �  CQ  	%�  F�,  	�u  H�,  	z  I�,  	ʓ  C�  ^  �>  =    	��  b�>  �   �>  =    	��  c�>  	0K  d�   	?�  e�   �	"?  x �Q   y �Q  dx �Q  dy �Q   ��  ��>  �P?  �p �
�.  ��  �
%1   �	?  {q �Q   ��  ��  d �	.?   t�  �P?  ?  �?  =   � 	r ��?  	�T  ��?  ?  	l�  �Q  	�  �Q  	?k  �Q  	�d  �Q  	2~ �"?  	��  ��  	��  �Q  	k�  �Q  	Z�  �%1  %1  5@  =    	�v  �%@  	�v  ��   	"�  ��.  �  �,  �U  {2  ��  {2  t�  �   �  	�   .Y  
Q  7Y  Q  �h  �@  �.  *� �.  <i  �.  	G  �  	��  �   �   	A  =    
K   �*A  )top  �G  �  �]  �	A   �	�A  ��  �%1   ��  �*A  O{  �
�   ��  �
�   iK  ��A   .  ��  �6A  �A  �A  =    	��  ��A  !K   �A  )up  �  �F  �S   FT  
�A  !K   B  ��   �x  H�  ��  �H   ��  �A  H	�B  `e �   >} <0  L� Q   $low Q  $+�  Q  (�Z !
�   ,r� "
�   0�f  #�A  4�f  $�A  8��  %�  <$tag &
�   @*� 'B  D �w )B  �B  �B  =    �B  �  2�B  !K   FAC  �c  +c �c d d �c hc �c  �c PC  @T	�C  `e V�   *� WAC  >} X<0   �}  YQ  (L� ZQ  ,��  ]�   0�c `�   4�c c�   8 �y eNC  !K   �
D  ��   �s  z�  ��  �T  ܭ   gY  ��C  H�	�D  `e ��   *� �
D  >} �<0   �W  �Q  (�}  �Q  ,L� �Q  0��  ��  4��  �
�   8$tag �
�   <��  �
�   @  w �D  �D  �D  =    �D  j�  �D  !K   X�D  )ok  �b �b  Mb ]�D  ) E  J @�E  � "�    � '
�@  �� *	�   
 -�E  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 E   H	�E  � K�    C� N	�   "8 QR   t TR    . V�E  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   E  KF    	R  @F  �E  bF    	�  WF  
K    rI  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	 !V�   ;6  	��  "M�  	(h  "N�   	l�  "N�   	�  #.�  	�  #/�  	�  #0�  	�  #2�  	w�  #8_  	�  #9&  	�  #:�  	�_  #;�   	��  #>�  	�  #J�  	"�  #R  	t�  #S�   	�w  #T�   	؜  #Y�   	q�  #[�  	Ƚ  #^  	�  #_�   	�y  #`�   	b�  #c�   	+�  #f�  	��  #i�  	֘ #l�   	�J  #x�   	��  #y�   	ks  #�   	�  #��   	J�  #��   	�i  #��   	��  #��  	��  #��  	��  #��  	<� #��  	��  #��  	��  #��  	5�  #��  	<m  #��   	 K  #��   	�R  #��   	op  #��   	�m  #��   	D  #��   	X�  #��   	If  #��   	� #��   	��  #��  	�U  #��  	`  #��  	J�  #��  	��  #��  	� #�@  �6  �K  =    	�  #��K  �  �K  =    	� #��K  ^  �K  =   	 	,�  #��K  	R�  #��K  ^  ^  L  =    	�u  #�L  	��  #��7  	�e  #��   �   JL  =   � 	(�  #�9L  	�  #��  ��  #@  �v  #�   n�  #�   4�  #�   *b #�   ��  #I  	Y�  $%�#  	��  $&�#  *�c }�@     n       �uM  +sec <0  �+ �+ ,�k  �   H, D, -Tw "uM  �, �, .��@     R  HM  /U@/T6/Q0 .��@     R  `M  /Us  0��@     )R  /Uv   �C  *"d +�@     R       ��M  +sec &<0  �, �, -Tw 	uM  - - .B�@     R  �M  /U@/T6/Q0 0M�@     R  /Us   *�c Q	�@     "      �TO  ,��  R%1  �- w- ,�p S�.  9. 5. -�R  U�9  z. r. 1sec V<0  �. �. -Tw WuM  / �. 2<p X
�    3�@            �N  -+w ��B  L/ J/  4��@     5R  �N  /U0/T" .7�@     AR  �N  /U	��B      5g�@     5R  .x�@     R  'O  /U@/T6/Q0 .��@     R  ?O  /Us  0�@     )R  /Uv   6�c ��   ڿ@     u      ��P  7��  �%1  u/ o/ 7*� �AC  �/ �/ -�k  
�   0 0 1rtn  �   �0 �0 1sec <0   1 1 -Tw uM  G1 C1 .�@     LR  P  /U~ /T|  .7�@     R  2P  /U@/T6/Q0 .B�@     R  JP  /Us  .��@     )R  bP  /Uv  .��@     )R  zP  /Uv  .��@     )R  �P  /Uv  .�@     )R  �P  /Uv  57�@     5R   67d ��   O�@     �       �SQ  7��  �%1  �1 }1 7*� �AC  2 �1 7�p ��.  �2 {2 8p ��9  �2 �2 .��@     5R  EQ  /U0/T" 9�@     TO   :vc 9)�@     �      �R  7Tw 9 uM  O3 33 8res ;�D  �4 {4 9��@     5R  .��@     XR  �Q  /R0/X1 .(�@     eR  �Q  /Us  .��@     XR  �Q  /R0/X1/Y1 ;׿@     eR  /U�U  <� � 6<3b 3b G<Ic Ic \	<� � !6=�E �E % <Vb Vb `>c c `<c c H R   =[  S#  j �*  ��@     �      k+ �m  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  9�  0t  4  e2    �0  }  ��  (  
K   J�  D   �C  
D  ���� �C  N\  ڵ  RP  �   	)  ��  "B   E�  #B  e% $I  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�  ;  
K   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (<  
K   /�  ��   [r  �4 #�  �   �X  5�  
K   :/  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K�  
�   Pn  =_  ��   R�  N�  ��  ��   �p  W;  
K   	3�  ��   ({  ��  ğ   F]  	8z  
K   	Y�  ��   �c  |  ��  l  ��  �   
K   	k7  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  	{�  
K   	�v  &�   �  º  GY  �f  ��   v�  	�C  
K   	��  GQ   ϼ  �  �_  X  &�  �b   t�  
 �   �  �  �  =   �' �  	��  1�  	]  4�  �  �    =   �    	Zy  8  �  8  =   =   � "  	��  ;8  Ʃ  QK   I  U  k  =     Z  	�  Wk  �p  #�  �  �   S�  $�  �  �  R    T}  %�  �  �  R   R    '	  acv )|  ��  *�  ��  +�   �y -�  �Y  6  ��  :O  s�  <O   �H  =O  xz  >     x @  I  q  =    ;  �  =    
�	�  x �I   y �I  Mp �I  *� �I  ޽  �I   ~x ��  
K   %
  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  
K   ��#  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u1
  (x	2$  �u z%
   � {	�   s |	�   � ~  N�  �#  ��  �	�   ��  �	�     J]  ��#  2$  P$  =   �  �^  �?$  �   h$  !  �  �]$  "K   ��'  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  u$  \	)  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /�'  )  8)  =   �  ��  1()  
K   p%*  �! 9& +! v( %# 0  B& @�! ��"  w#  	$  �-  S%  �)   0  @&  ��"    !0    m0    b-    �.    �$     /   @ %   � <"    U-    5'    	!  �]  ���+  `e �U   x ��  y ��  z ��   ��  ��+  (cN  ��+  0Mp �I  8�u �%
  <� ��   @�H  ��+  Hr�  ��+  P��  �6,  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� ��'  �y� �<,  �s ��   ��� �B,  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  �+  ���  �   ���  	�   ��R  ".  �f�  �   �I}  �  ���  �+  � %*  Gx  �6,  >} ��1   �}  �I  �|  �I  
 ,  )  2$  #d  HN".  mo P@0   ��  Q;7  cmd R)  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  gG7  8�W  hW7  P��  i�  h�� lF0  l�N  m7  |E�  p7  ��W  rg7  �~�  sF0  �*� tF0  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �@0  �$�R  ��    $��  ��   $�  ��   $h  �w7  $I�  ��  @ H,  �z %*  �  	��  ��   	�\  ��  	�  �_.  �  	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  �5.  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	/  x E�   y F�   �{ H�.  (T	Z/  `e VU   x W�  y X�  z Y�    	�  ["/  �a	@0  = c�   F�  d�  �~ eI  h�  fI  
t�  gI  �k hI  tag iI  �N  l
�   ��  o@0  ��  r
F0   iK  uZ/  0��  x
�   XS�  {@0  `��  ~R   h��  ��   pu| �1  x (.  �   V0  =    �}  X�1  v1 ��1   v2 ��1  dx ��  dy ��  �  �I  �k �I  tag �I  �W  �a  �o ��1  $��  ��1  4SX  ��1  8d�  ��1  @��  �
�   H��  �R   P 1  V0  �z �f/  �	�1  2�  ��   ]  ��  �h  �I  �N  �I  
�K  �I  >} ��1   "1  �}  �.1  
K   ��1  ��   �  o�  ��   ��  ��1  /  �  �1  =    �u  �V0  �z �,  8�	i2  v1 ��1   v2 ��1  82  ��  Mp �I  [�  �i2   �  �o2   SX  ��1  (d�  ��1  0 �1  �1  A{ ��1  4	�2  %x �   %y 	�  %dx 
�  %dy �  �o �2  )�  q  0 �  �2  =   =    (} �2  �  *�  &v  @2�3  @�  4�3   %x1 5�   %x2 6�   .]  8�  5]  9�  �� :�  ��  =�   �  @�   ��  C�  $�n  G�3  (9x  H�3  0�^  I�3  8 u2  I  >�  K
3  &�h  PR�4  s�  U�4   �H  V�4  %x1 X�   %x2 Y�   %gx \�  %gy ]�  %gz `�   %gzt a�  $�x  d�  (� f�  ,~�  i�  0t  k�  4.� l�   8�  p�4  @	�  r�   H �3  �2  �h  t�3  �	5  �c  ��   �O  �5  �x  �
5   I  5  =    �  "5  =    I�  ��4  �	V5  �  ��    �  �V5   "5  �  �/5  '��	6    ��   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  %top �	6  (��  �	�  U(��  �	�  V(� �	6  W(�  �	�  � �  $6  =   ? ��  �i5  	�6  ~�  v   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %16  �6  �6  =    	S�  '�6  
K   7�6  {�   U�  ~�   >	7  �� @B,   s A
�   sx B�  sy C�   Nz E�6  
K   1;7  ��   ��  ��   �y  97  �   W7  =    �  g7  =    �  w7  =    7  �7  =    hy �H,  (�	�7  in ��   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
F0  �a  �
�   $ ��  ��7  ��	�8  2�  �
�    I�  ��  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��8  ( �7  �8  =    ޴  �8  	.L  &�8  �  	׮  )�8  	�  +�8  	�  ,�8  	�Q  .�4  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  769  �   	��  869  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�9  \5  	��  H�   	��  I�1  	��  K�   	a� L�3  	w�  N�   	P{ O�1  	��  Q�   	��  R�9  �1  	��  T�   	�� U:  �2  	�}  W�   	u| Xo2  	M�  Z�   	P�  [i2  	��  a�  	��  b�  	�  c�  	�p  eI  	�T  fz:  �7  	�a  jI  �   �:  =   � 	ը  l�:  I  �:  =   @ 	�p  m�:  	 �  p�  	p|  qI  	$Y  v�   	�K  y�   	g  {;  $6  	d�  |;  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   �4  �;  =   =   / 	��  E�;  �4  �;  =   / 	Ԁ  F�;  �4  �;  =   =    	7� G�;  	�R  I�   	��  J�4  	��  U�   	P�  \5  	��  ]5  	L�  ^5  	ߵ  _5  	�  a5  	@�  �3  	[�  i2  	 �  o2  	SX  �1  	d�  �1  	��  �   	_�   �   	��  "�  	��  %�  	'�  &�  	�]  (�  �3  �<  =   � 	�P  *�<  	ӯ  +=  �3  	|  -"=  �4  	��  ."=  	��  /"=  F=  V=  �   �    	��  �3  �   @=  	qY  "b=  	�  #b=  I  �=  =   ? 	��  %�=  	��  &�=  �  �=  =   � 	@Y  (�=  �  �=  =   ? 	V�  )�=  �4  �=  =    	�h  �=  	�  >  �4  	�  �4  	�f  !�=  	r�  "�=  	��  %�3  	��  &�3  	׆  '�  	��  (�  	�  *�  	��  +�  	�  �4  	��  �   	�_  �   	�_  �   	b  �  	t  �  	j�  "5.  	�  :�   	��  ;�   	��  <�   	�W  >�4  	hn  @�  	U~  A�  	�  B�  	 �  C�  	%�  F5.  	�u  H5.  	z  I5.  	ʓ  CU  �  v?  =    	��  bf?  �   �?  =    	��  c�?  	0K  d�   	?�  e�   �	�?  x ��   y ��  dx ��  dy ��   ��  ��?  �@  �p �
@0  ��  �
o2   �	K@  {q ��   ��  ��  d �	�?   t�  �@  K@  g@  =   � 	r �W@  	�T  �@  K@  	l�  ��  	�  ��  	?k  ��  	�d  ��  	2~ ��?  	��  ��  	��  ��  	k�  ��  	Z�  �o2  o2  A  =    	�v  ��@  	�v  ��   	"�  �@0   �  5.   �U  �3   ��  �3   t�  �    �  	�    .Y  
�   7Y  �   �h  �A  @0   *� F0   <i  F0  	G  �  	��  �   �   �A  =    
K   ��A  )top  �G  �  �]  ��A   �	MB  ��  �o2   ��  ��A  O{  �
�   ��  �
�   iK  �MB   Z/  ��  �B  SB  oB  =    	��  �_B  "K   �B  )up  �  �F  �S   FT  
{B  "K   �B  ��   �x  H�  ��  �H   ��  �B  H	�C  `e U   >} �1  L� �   %low �  $+�  �  (�Z !
�   ,r� "
�   0�f  #�B  4�f  $�B  8��  %�  <%tag &
�   @*� '�B  D �w )�B  �C  �C  =    �C   �  2�C  "K   FD  �c  +c �c d d �c hc �c  "K   �AD  ��   �s  z�  ��  �T  ܭ   gY  �D  H�	�D  `e �U   *� �AD  >} ��1   �W  ��  (�}  ��  ,L� ��  0��  ��  4��  �
�   8%tag �
�   <��  �
�   @  w �ND  E  E  =    �D   j�  �D  "K   sE  �g  Fe 	h g qf �j �e �f �h i 	�j 
�h ]h  ) E  J @F  � "�    � '
�A  �� *	�   
 -F  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 sE   H	SF  � K�    C� N	�   "8 QR   t TR    . VF  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   sE  �F  ! 	R �F  SF  �F  ! 	� �F  
K   rxI  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	 V�   	�  M�   	5  N�   )  	��  !M�  	(h  !N�   	l�  !N�   	�  ".�  	�  "/�  	�  "0�  	�  "2�  	w�  "8�  	�  "9�  	�  ":/  	�_  ";�   	��  ">�  	�  "J�  	"�  "Rn  	t�  "S�   	�w  "T�   	؜  "Y�   	q�  "[�  	Ƚ  "^n  	�  "_�   	�y  "`�   	b�  "c�   	+�  "f�  	��  "i�  	֘ "l�   	�J  "x�   	��  "y�   	ks  "�   	�  "��   	J�  "��   	�i  "��   	��  "��  	��  "��  	��  "��  	<� "��  	��  "��  	��  "��  	5�  "��  	<m  "��   	 K  "��   	�R  "��   	op  "��   	�m  "��   	D  "��   	X�  "��   	If  "��   	� "��   	��  "��  	�U  "��  	`  "��  	J�  "��  	��  "��  	� "��  �7  .L  =    	�  "�L  �  JL  =    	� "�:L  �  fL  =   	 	,�  "�VL  	R�  "�~L  �  �  �L  =    	�u  "��L  	��  "��8  	�e  "��   �   �L  =   � 	(�  "��L  	�  "��   ��  "�   �v  "�    n�  "�    4�  "�    *b "�    ��  "�I  
K   -zM  �g  �g sg Ih �h �f �i he �h �e 	 1e 9/M  zM  �M  =    *k ?�M  	@[e     zM  �M  =    *�j E�M  	 [e     *��  `
@0  	8Hf     �  �M  =    +�d 	�M  	 [e     +~j 	�M  	�Ze     +;e ��   	�Ze     +zd U
@0  	(Hf     +h V
@0  	0Hf     +�j W
�  	@Hf     +�g X
�  	DHf     @0  �N  =    +h 
�N  	`Hf     +h �   	 Hf     +�d �   	�e     ,Ud �h�@     #       �DO  -mo �@0  �4 �4 .*u �
�   5 5 /��@     �}   0j ��O  1mo �@0  20g �@0  3fog �@0  2:J �@0  3r �
�   2*� ��'   ,�i �Q�@            �P  -mo �@0  K5 C5 4_�@     �}  �O  5Us 5T_ 6h�@     DO  5U�U  ,�g k��@     �       ��P  -mo k@0  �5 �5 .:J m@0  6 6 .0g n@0  Q6 M6 7U�  p�   	�e     4�@     ~  �P  5Us 5Tv 5QL 6H�@     �}  5U05T^  ,�i f��@            ��P  -mo f@0  �6 �6 /��@     ~   ,�j Q=�@     �       ��Q  -mo Q@0  �6 �6 8x S
�   7 7 8y T
�   ?7 ;7 8z U
�   y7 u7 8th V@0  �7 �7 9M�@     ~  9T�@     ~  9^�@     ~  4{�@     %~  �Q  5Us 5Tv 5R! 9��@     ~  4��@     1~  �Q  5Us 5T
 9��@     ~   ,�f 7��@     �       � S  -mo 7@0  �7 �7 8x 9
�   D8 B8 8y :
�   i8 g8 8z ;
�   �8 �8 8th <@0  �8 �8 9��@     ~  4��@     %~  �R  5Us 5T| 5R! 9��@     ~  4�@     1~  �R  5U| 5T
 9�@     ~  6=�@     �}  5U05Tb  ,nd 1��@            �MS  -mo 1@0  9 9 6��@     �}  5U05Ta  ,�f &�@     e       ��S  -mo @0  H9 D9 .`e �S  �9 �9 8m @0  �9 �9 6��@     �}  5U05T`  U  ,kh �@     $       �ET  :�R  z:  �9 �9 -psp ET  :: 2: 4�@     �}  (T  5T6 6&�@     =~  5U�U5T�T  7  ,!g ���@            ��T  :�R  �z:  �: �: -psp �ET  �: �: 6�@     �}  5T7  ,{h ���@            �U  :�R  �z:  ; ; -psp �ET  T; P; 6��@     �}  5T5  ,e ���@            �lU  -mo �@0  �; �; 4��@     �}  VU  5Us 5TO 6��@     0o  5U�U  ,�i ���@            ��U  -mo �@0  �; �; 4��@     �}  �U  5Us 5TU 6��@     0o  5U�U  ,4i ���@            �:V  -mo �@0  c< [< 4��@     �}  $V  5Us 5TT 6��@     0o  5U�U  ,j x��@     �      �'W  -mo x@0  �< �< 8th z�S  r= n= 8mo2 {@0  �= �= 7,e |�1  ��8i }
�   �= �= ;'W  9�@      �  ��V  <9W  "> >  4~�@     J~  �V  5U�� 4��@     W~  W  5U��5T6 9��@     ~   =�e E�  GW  >�j E(�'   ,$h :��@            ��W  :�g :@0  \> X> 6��@     d~  5U�U5Q�  0�h -�W  >�d -@0   ,Ui %��@            ��W  :�d %@0  �> �> 6��@     �}  5U�U  ,e  ��@     
       �LX  :�d  @0  �> �> 6��@     �}  5U�U5TO  ,�d �g�@     `       ��X  :�d �@0  .? $? .*u �
�   �? �? 9��@     ~  9��@     ~  /��@     �}   ,
f �+�@     <       �_Y  :�d �@0  �? �? ;�W  +�@     �  �Y  <�W  C@ A@  4D�@     �Y  1Y  5Us  4U�@     �Y  IY  5Us  6g�@     �Y  5U�U  ,�i ��@             ��Y  :�d �@0  p@ f@ 4�@     o  �Y  5Us  6*�@     �Y  5U�U  0�h �KZ  >�d �@0  >Mp �I  3x ��  3y ��  3z ��  20g �@0  3an �I  2=f �
�   2r� �
�   2Ye ��S   ,0j �`�@     �       �-[  :�d �@0  �@ �@ .`5 �@0  6A 4A 8an �I  [A YA .S� ��   �A ~A 4��@     �}  �Z  5Us  4��@     o  �Z  5Us  4��@     p~  [  5UD@$ 4��@     p~  [  5UD@$ 9��@     |~   ,�e i��@     �       �>\  :�d i@0  �A �A 8mo k@0  BB :B . �  l@0  �B �B 8an m
�   �B �B 4��@     o  �[  5U|  9��@     �~  4��@     ~  �[  5U| 5T} 5Q9 9��@     p~  9��@     p~  4�@     ~  #\  5U| 5T} 5Q9 9<�@     p~  9U�@     p~   ,�e V��@     �       �5]  :�d V@0  C C 8mo X@0  hC dC . �  Y@0  �C �C 8an Z
�   �C �C 4��@     o  �\  5Us  9�@     �~  4!�@     ~  �\  5Us 5Tv 5Q9 41�@     ~  ]  5Us 5Tv 5Q9 9a�@     p~  9z�@     p~   ,�e B_�@     �       �,^  :�d B@0  D �C 8mo D@0  SD OD . �  E@0  �D �D 8an F
�   �D �D 4j�@     o  �]  5Us  9}�@     �~  4��@     ~  �]  5Us 5Tv 5Q9 4��@     ~  ^  5Us 5Tv 5Q9 9��@     p~  9��@     p~   ,Ji ;H�@            ��^  :�d ;@0  �D �D 4Q�@     o  x^  5Us  6_�@     �}  5U�U5Tc  ,Dg [�@     �       ��_  :�d @0  ]E OE .��  @0  �E �E 8an 
�   4F 2F 4x�@     o  	_  5Us  4��@     �~  !_  5Us  4��@     �}  ?_  5Us 5TR 4��@     �~  b_  5Ts 5Qs 5RD 4��@     p~  {_  5UH@$ 4 �@     p~  �_  5UH@$ 6?�@     d~  5T�U5QF  ,�d �	�@     R       �6`  :�d �@0  gF ]F 8fog �@0  �F �F 4�@     o  `  5Us  45�@     %~  (`  5R4 /Z�@     6`   ,�g �A�@     �       �-a  :�d �@0  G  G .`5 �@0  kG gG . �  �@0  �G �G 8an �K   �G �G 9c�@     �~  4n�@     �~  �`  5Tv  4~�@     �~  �`  5Us  4��@     p~  �`  5UH@$ 4��@     p~  a  5UH@$ 6��@     �~  5U�U  ,�g ���@            ��a  :�d �@0  �G �G 4 �@     �}  a  5Us 5T[ 6	�@     6`  5U�U  ,=h ���@            ��a  :�d �@0  ZH RH 4��@     �}  �a  5Us 5T\ 6��@     6`  5U�U  ,�f �7�@     
       �Mb  :�d �@0  �H �H 6A�@     �}  5U�U5T6  ,�f ���@     e      ��c  :�d �@0  I �H 8xl ��   �I �I 8xh ��   �I �I 8yl ��   �I �I 8yh ��   'J #J 8bx ��   aJ ]J 8by ��   �J �J .y� �<,  �J �J .v� �@0  �J �J 4��@     �~  Nc  5U~ 5T 5Q	��@      4��@     o  fc  5Uv  4��@     1~  �c  5Uv 5T

 4��@     �}  �c  5TO 9��@     1~  67�@     0o  5U�U  ?�d Z	�  �c  >�p Z @0  2�i \
�   2Wy ]�   ,�f >j�@     h       ��d  :�d >@0  )K K .\q @
�   �K �K 4��@     o  Zd  5Us  4��@     �u  rd  5Us  9��@     ~  4��@     �}  �d  5Us 5T5 6��@     �~  5T�U5Q�U5R�l�:#6  ,�j 6H�@     "       �4e  :�d 6@0  "L L 4[�@     o  e  5Us  6i�@     �}  5U�U5T8  ,�e ���@     `      �6f  :�d �@0  �L �L .�f �I  �L �L .S� ��  9M 5M .�  ��  �M �M .`5 �@0  �M �M 8th �@0  �M �M 9
�@     �~  4#�@     %~  �e  5R7 92�@     ~  9}�@     �~  9��@     p~  9��@     p~  9�@     |~   ,�d ���@     R       ��f  :�d �@0  -N %N 8mo �@0  �N �N 4��@     o  �f  5Us  @��@     ~  5Us 5Q6  ,!f �7�@     _       �wg  :�d �@0  �N �N .\q �
�   sO oO 4J�@     �u  g  5Us  4[�@     �}  /g  5Us 5T7 9`�@     ~  A��@     �~  \g  5T�U5Q�U 6��@     ~  5U�U5Q@  ,�i ��@     )       ��g  :�d �@0  �O �O 4!�@     o  �g  5Us  66�@     ~  5U�U5Q!  ,�i ���@     Z       ��h  :�d �@0  AP 1P .\q �
�   �P �P 4��@     o  @h  5Us  4��@     �u  Xh  5Us  9��@     ~  A��@     �~  �h  5T�U5Q�U 6�@     ~  5U�U5Q   ,fi �k�@     I       �Di  :�d �@0  CQ 5Q .\q �
�   �Q �Q 4~�@     o  i  5Us  4��@     �u  i  5Us  9��@     ~  6��@     �~  5T�U5Q�U  ,/f ��@     g       �#j  :�d �@0  R R .\q �
�   �R �R 4�@     o  �i  5Us  4�@     �u  �i  5Us  40�@     �}  �i  5Us 5T7 95�@     ~  AU�@     �~  j  5T�U5Q�U 6j�@     ~  5U�U5QO  ,�g s��@     )       ��j  :�d s@0  S �R 4��@     o  oj  5Us  6�@     ~  5U�U5Q$  ,�d c��@     I       �k  :�d c@0  �S zS 4��@     o  �j  5Us  9��@     ~  A��@     1~  �j  5U�U @��@     �~  5Us   ,�i RI�@     I       ��k  :�d R@0  T T 4R�@     o  ^k  5Us  9W�@     ~  A{�@     1~  �k  5U�U @��@     �~  5Us   ,	g >��@            ��l  :�d >@0  �T �T .Mp @
�   "U U .|e A
�   ZU XU .\q B
�   U }U .�  C
�   �U �U 4��@     �}  >l  5Us 5T2 4��@     o  Vl  5Us  4�@     �~  {l  5Us 5T} 5Q@G$ 9�@     ~  9�@     ~  9�@     ~  6H�@     �~  5U�U5Q@G$  ,qj &2�@     �       �n  :�d &@0  V �U 8i (
�   jV dV .Mp )
�   �V �V .|e *
�   �V �V .\q +
�   W 	W .�  ,
�   >W :W 4d�@     �}  wm  5Us 5T2 4l�@     o  �m  5Us  4��@     �~  �m  5Us 5T} 5Q@G$ 9��@     ~  9��@     ~  9��@     ~  @��@     �~  5Us 5Tv 5Q@G$5R~   ,i ��@            �o  :�d @0  ~W tW .Mp 
�   �W �W .\q 
�   AX ?X .�  
�   vX pX 4��@     o  �n  5Us  4��@     �~  �n  5Us 5T} 5Q@G$ 4��@     �}  �n  5Us 5T1 9��@     ~  9��@     ~  9�@     ~  61�@     �~  5U�U5Q@G$  0#j �0o  >�d �@0   ,�e �f�@     �      ��p  :�d �@0  �X �X .� �
�   �Y �Y B�g ���@     4��@     ir  �o  5Us 5T1 AD�@     Gs  �o  5U�U 4Y�@     �u  �o  5Us  4s�@     �}  �o  5Us  A��@     1~  	p  5U�U 4��@     eu  !p  5Us  4��@     1~  9p  5Us  4�@     �~  Qp  5Us  4�@     ir  np  5Us 5T1 4%�@     u  �p  5Us  41�@     Gs  �p  5Us  9C�@     ~  6[�@     �}  5U�U  ,�i M��@     �       ��q  :�d M@0  Z �Y .:J O@0  �Z �Z BVh g��@     C�@     I       mq  .*u j�   �Z �Z 9�@     ~  9.�@     ~  9Q�@     �}   4��@     ir  �q  5Us 5T0 9�@     �~  6d�@     1~  5U�U  ,dd 'A�@     b       �ir  -mo '@0  [ [ 8th )�S  o[ k[ 8mo2 *@0  �[ �[ 7,e +�1  ��D�W  A�@     A�@            -Nr  <�W  �[ �[  @��@     W~  5U��5T3  E`f ��  )�@           �Gs  :�d �@0  
\ \ :�g ��  \\ V\ 8c �
�   �\ �\ .�� �
�   $] "] 2�R  �z:  8an �I  K] I] .S� ��  w] u] 4��@     �~  ,s  5Us  9��@     �~  9�@     |~   ,>j _��@     D      ��t  :�d _@0  �] �] .Gd a�  �] �] .Nd b�  ~^ z^ 8d d�t  �^ �^ .�j f
�   �_ �_ .�d gzM  �_ �_ .Lj izM  #` !` 4�@       t  5U	�B      4��@     �t  .t  5Us  9��@     ~  4 �@     �t  St  5Us  4F�@     �t  kt  5Us  4a�@     �t  �t  5Us  9n�@     ~  4��@     �t  �t  5Us  4��@     �t  �t  5Us  @��@     �t  5Us   zM  �t  =    ?"e Q	�  u  >�d Q@0   ?ue 	�  eu  >�d @0  2�j �  2�g �  3ld 	o2  2�j �  2|g �   F�d �	�  �u  G�d �&@0  HS� ��   FQg �	�  �u  G�d �$@0  Ipl �@0  HS� ��   JWj �3�@            �v  K �  �@0  L` F` K�j �@0  �` �` 6N�@     v  5T0  Lsi cfv  Msec d�1  G8g e�   Ii g
�   HWy ho2  H�  i�1   N�c  ��@     �       ��v  <�c  �` �` O�c  O�c  P�c  �  <�c  3a /a Q�  R�c  na la R�c  �a �a @m�@       5U�U    Nv  ��@     �       ��w  <+v  �a �a <7v  %b b RCv  �b �b OMv  OYv  Sv  ��@     p       <7v  �b �b <+v  �b �b T��@     p       RCv  *c $c RMv  wc uc RYv  �c �c 4��@       �w  5U|  9%�@     v     N�u  N�@     V       �gx  <�u  �c �c R�u  @d >d R�u  ed cd U�u  ��@            Yx  <�u  �d �d T��@            O�u  O�u  @��@     �~  5Us    9u�@     |~   Neu  ��@           �	y  <vu  �d �d O�u  Ueu  ��@     �       �x  <vu  e �d T��@     �       R�u  4e $e 9��@     |~  9��@     ~    @��@     �~  5Uv   Nu  ��@           �	z  <u  �e �e R$u  ff bf R1u  �f �f O>u  RJu  ng fg OWu  Uu  �@     �       �y  <u  �g �g T�@     �       O$u  O1u  O>u  OJu  RWu  �g �g @��@     %  5Us 5Q0   4��@       �y  5U	��B      @�@     1  5Us   N�t  ��@     "       �zz  <�t  0h *h U�t  ��@            ez  <�t  ~h |h 9��@     ~   @��@     u  5Us   No  ]�@     V       ��z  <"o  �h �h Uo  ��@            �z  <"o  
i i 9��@     ~  9��@     ~   9��@     �~   N�Y  �@     �       �z|  <�Y  ;i -i <�Y  �i �i O�Y  O�Y  O�Y  O
Z  OZ  O#Z  R0Z  .j (j R=Z  |j xj P�Y  0  <�Y  �j �j <�Y  k k Q0  R�Y  �k �k R�Y  �k �k R�Y   l �k R
Z  Hl >l RZ  �l �l R#Z  'm %m O0Z  O=Z  4��@     p~  �{  5Us  4��@     p~  |  5Us  4��@     %~  +|  5U} 5RB 4��@     1  C|  5Us  A��@     �~  j|  5T�U5Q�U5R
' /
�@     KZ     N�W  ��@            ��|  V�W  U NDO  I�@           ��}  <RO  Tm Jm O^O  OkO  OxO  O�O  O�O  PDO     <RO  �m �m Q   R^O  1n -n RkO  in gn RxO  �n �n R�O  �n �n R�O  �n �n 9g�@     �~  4}�@     %~  ^}  5RM 4��@     �}  v}  5T# 9��@     ~  9�@     %~  4!�@     ir  �}  5Us 5T1 47�@     1~  �}  5Us  4E�@     =  �}  5Us  6P�@     I  5U�U    W� � 6W�j �j x	W�. �.  <W� � #!W�( �( kW�e �e s	X�h �h  XUf Uf nX�c �c rW.h .h �Wd  d  
"	W�h �h �	W�e �e r	W�f �f �	Xdj dj Wi i �W�d �d �W�h �h �	W�e �e vWEf Ef xWcg cg �Wf f �W��  ��  $7W�" �" �	W�g �g �W�i �i 1W\i \i �	W;i ;i �	W11 11 q ,T   X`  S#  �k �*  ��@     �      �J �p  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  
K   "f  ��  WH  �~  �O  �m  ��   �  ��  ��  	 0t  r  e2    �0  }  ��  f  
K   J�  D   �C  
D  ���� �C  N�  ڵ  R�  �  
K   &  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
K   /_  ��   [r  �4 #�  �   �X  52  
K   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  Kk  
�   P  =_  ��   R�  N�  ��  ��   �p  W�  
K   	3@  ��   ({  ��  ğ   F]  	8  
K   	k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  	{L  
K   	��  &�   �  º  GY  �f  ��   v�  	��  t�  
 �   �  �  
  =   �' �  	��  1
  	]  4'  �  �  >  =   � -  	Zy  8>  �  e  =   =   � O  	��  ;e  Ʃ  QK   v  �  �  =     �  	�  W�  �p  #�  �  �   S�  $�  �  �  R    T}  %�  �    R   R    '	/  acv )�  ��  *�  ��  +�   �y -  �Y  6/  ��  :|  s�  <|   �H  =|  xz  >;   G  x @G  �  �  =    y  �  =    
�	�  x ��   y ��  Mp ��  *� ��  ޽  ��   ~x ��  
K   R	  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �  
K   ��"  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u^	  (x	_#  �u zR	   � {	�   s |	�   � ~/  N�  �"  ��  �	�   ��  �	�     J]  ��"  _#  }#  =   � �^  �l#  �   �#    �  ��#  !K   ��&  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �#  \	H(  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /�&  H(  e(  =   � ��  1U(  �]  ��H*  `e ��   x ��  y ��  z ��   ��  �H*  (cN  �H*  0Mp �v  8�u �R	  <� ��   @�H  �H*  Hr�  �H*  P��  ��*  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� ��&  �y� ��*  �s ��   ��� ��*  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  H*  ���  �   ���  	�   ��R  o,  �f�  �   �I}  �  ���  H*  � r(  Gx  ��*  >} ��/   �}  ��  �|  ��  
 N*  H(  _#  "d  HNo,  mo P�.   ��  Q�5  cmd R�5  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g6  8�W  h6  P��  i�  h�� l�.  l�N  m�  |E�  p�  ��W  r+6  �~�  s�.  �*� t�.  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��.  �#�R  ��    #��  ��   #�  ��   #h  �;6  #I�  ��  @ �*  �z r(  �  	��  ��   	�\  ��  	�  ��,  �  	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  ��,  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	c-  x E�   y F�   �{ HC-  (T	�-  `e V�   x W�  y X�  z Y�    	�  [o-  �a	�.  = c�   F�  d�  �~ e�  h�  f�  
t�  g�  �k h�  tag i�  �N  l
�   ��  o�.  ��  r
�.   iK  u�-  0��  x
�   XS�  {�.  `��  ~R   h��  ��   pu| �c/  x u,  �   �.  =    �}  X�c/  v1 �0   v2 �0  dx ��  dy ��  �  ��  �k ��  tag ��  �W  ��  �o �0  $��  �0  4SX  ��/  8d�  ��/  @��  �
�   H��  �R   P i/  �.  �z ��-  �	�/  2�  ��   ]  ��  �h  ��  �N  ��  
�K  ��  >} ��/   o/  �}  �{/  
K   �0  ��   �  o�  ��   ��  ��/  c-  �  .0  =    �u  ��.  �z �N*  8�	�0  v1 �0   v2 �0  82  ��  Mp �v  [�  ��0   �  ��0   SX  ��/  (d�  ��/  0 �/  .0  A{ �F0  4	'1  $x �   $y 	�  $dx 
�  $dy �  �o '1  )�  �  0 �  =1  =   =    (} �0  �  *�  %v  @22  @�  42   $x1 5�   $x2 6�   .]  8�  5]  9�  �� :�  ��  =�   �  @�   ��  C�  $�n  G2  (9x  H2  0�^  I2  8 �0  �  >�  KW1  %�h  PR3  s�  U3   �H  V3  $x1 X�   $x2 Y�   $gx \�  $gy ]�  $gz `�   $gzt a�  $�x  d�  (� f�  ,~�  i�  0t  k�  4.� l�   8�  p3  @	�  r�   H %2  J1  �h  t%2  �	O3  �c  ��   �O  �O3  �x  �
_3   �  _3  =    �  o3  =    I�  �3  �	�3  �  ��    �  ��3   o3  �  �|3  &��	`4    ��   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  $top �	`4  '��  �	�  U'��  �	�  V'� �	`4  W'�  �	�  � �  q4  =   ? ��  ��3  	�4  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %~4  �4  �4  =    	S�  '�4  >	:5  �� @�*   s A
�   sx B�  sy C�   Nz E�4   	�5  ��  "�   E�  #�  e% $�  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4F5  
K   1�5  ��   ��  ��   �y  9�5  �   6  =    �  +6  =    �  ;6  =    :5  K6  =    hy ��*  (�	�6  in ��   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�.  �a  �
�   $ ��  �W6  ��	`7  2�  �
�    I�  ��  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  �`7  ( �6  p7  =    ޴  ��6  	.L  &�7  �  	׮  )�7  	�  +�7  	�  ,�7  	�Q  .3  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�7  �   	��  8�7  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u FH8  �3  	��  H�   	��  I0  	��  K�   	a� L2  	w�  N�   	P{ O�/  	��  Q�   	��  R�8  :0  	��  T�   	�� U�8  =1  	�}  W�   	u| X�0  	M�  Z�   	P�  [�0  	��  a�  	��  b�  	�  c�  	�p  ev  	�T  f>9  K6  	�a  jv  �   a9  =   � 	ը  lP9  v  ~9  =   @ 	�p  mm9  	 �  p�  	p|  qv  	$Y  v�   	�K  y�   	g  {�9  q4  	d�  |�9  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   3  ~:  =   =   / 	��  Eh:  3  �:  =   / 	Ԁ  F�:  3  �:  =   =    	7� G�:  	�R  I�   	��  J3  	��  U�   (	P�  \�:  �:  	��  ]�:  	L�  ^�:  	ߵ  _�:  	�  a�:  	@�  2  	[�  �0  	 �  �0  	SX  �/  	d�  �/  	��  �   	_�   �   	��  "�  	��  %�  	'�  &�  	�]  (�  2  �;  =   � 	�P  *�;  	ӯ  +�;  2  	|  -�;  3  	��  .�;  	��  /�;  <  !<  �   �    	��  2  �   <  	qY  "-<  	�  #-<  �  b<  =   ? 	��  %Q<  	��  &Q<  �  �<  =   � 	@Y  (z<  �  �<  =   ? 	V�  )�<  3  �<  =    	�h  �<  	�  �<  3  	�  3  	�f  !Q<  	r�  "Q<  	��  %2  	��  &2  	׆  '�  	��  (�  	�  *�  	��  +�  	�  3  	��  �   	�_  �   	�_  �   	b  �  	t  �  	j�  "�,  	�  :�   	��  ;�   	��  <�   	�W  >3  	hn  @�  	U~  A�  	�  B�  	 �  C�  	%�  F�,  	�u  H�,  	z  I�,  	ʓ  C�  �  A>  =    	��  b1>  �   ]>  =    	��  cM>  	0K  d�   	?�  e�   �	�>  x ��   y ��  dx ��  dy ��   ��  ��>  ��>  �p �
�.  ��  �
�0   �	?  {q ��   ��  ��  d �	�>   t�  ��>  ?  2?  =   � 	r �"?  	�T  �J?  ?  	l�  ��  	�  ��  	?k  ��  	�d  ��  	2~ ��>  	��  ��  	��  ��  	k�  ��  	Z�  ��0  �0  �?  =    	�v  ��?  	�v  ��   	"�  ��.  �  �,  �U  2  ��  2  t�  �   �  	�   .Y  
�  7Y  �  �h  X@  �.  *� �.  <i  �.  	G  �  	��  �   �   �@  =    
K   ��@  )top  �G  �  �]  ��@   �	A  ��  ��0   ��  ��@  O{  �
�   ��  �
�   iK  �A   �-  ��  ��@  A  :A  =    	��  �*A  !K   mA  )up  �  �F  �S   FT  
FA  !K   �A  ��   �x  H�  ��  �H   ��  zA  H	hB  `e �   >} �/  L� �   $low �  $+�  �  (�Z !
�   ,r� "
�   0�f  #mA  4�f  $mA  8��  %�  <$tag &
�   @*� '�A  D �w )�A  �B  �B  =    hB  �  2uB  !K   ��B  ��   �s  z�  ��  �T  ܭ   gY  ��B  H�	pC  `e ��   *� ��B  >} ��/   �W  ��  (�}  ��  ,L� ��  0��  ��  4��  �
�   8$tag �
�   <��  �
�   @  w ��B  �C  �C  =    pC  j�  }C  !K   �C  �g  Fe 	h g qf �j �e �f �h i 	�j 
�h ]h  �k 7�C  !K   ='D  1l  �k  �k AD  @E	�D  `e G�   *� H�C  ��  I�  >} J�/   ��  K
�   (}k L
�   ,P{  M�  0l N�  4L� O�  8 �x Q4D  !K   X�D  )ok  �b �b  Mb ]�D  ) E  J @�E  � "�    � '
�@  �� *	�   
 -�E  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 �D   H	�E  � K�    C� N	�   "8 QR   t TR    . V�E  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   �D  7F    	R ,F  �E  NF    	� CF  
K   r�H  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	  V�   �5  	��  !M�  	(h  !N�   	l�  !N�   	�  ".�  	�  "/�  	�  "0�  	�  "2�  	w�  "8_  	�  "9&  	�  ":�  	�_  ";�   	��  ">�  	�  "J�  	"�  "R  	t�  "S�   	�w  "T�   	؜  "Y�   	q�  "[�  	Ƚ  "^  	�  "_�   	�y  "`�   	b�  "c�   	+�  "f�  	��  "i�  	֘ "l�   	�J  "x�   	��  "y�   	ks  "�   	�  "��   	J�  "��   	�i  "��   	��  "��  	��  "��  	��  "��  	<� "��  	��  "��  	��  "��  	5�  "��  	<m  "��   	 K  "��   	�R  "��   	op  "��   	�m  "��   	D  "��   	X�  "��   	If  "��   	� "��   	��  "��  	�U  "��  	`  "��  	J�  "��  	��  "��  	� "�@  K6  �K  =    	�  "��K  �  �K  =    	� "��K  �  �K  =   	 	,�  "��K  	R�  "��K  �  �  L  =    	�u  "��K  	��  "�p7  	�e  "��   �   6L  =   � 	(�  "�%L  	�  "��  ��  "@  �v  "�   n�  "�   4�  "�   *b "�   ��  "	I  *�k ��   �@     �      �rN  +��  ��0  o o +*� �'D  ho bo ,�k ��   �o �o ,  ��   �p �p -i ��   �p �p ,�k ��   Bq :q ,P{  ��   �q �q -ok ��   r �q -rtn ��   Wr Mr -sec ��/  �r �r ,�k ��/  Is Cs ,�v �rN  �s �s ,�k ��  t t ,L� ��  ht `t .��@     �S  N  /Uw /Tv  .��@     �S  #N  /U@/T6/Q0 .��@     �S  ;N  /U~  .��@     �S  ]N  /U@/T6/Q0 0��@     �S  /Us   �D  1Uf ��   (�@     W      �Q  2��  ��0  �t �t 2-k ��C  u u 3�k ��   uu iu -rtn  �   v �u -i �   xv tv -sec �/  �v �v ,�v rN  w w 4@�@     �       �O  ,7k m�   Pw Lw ,<p n�0  �w �w .k�@     �S  �O  /Us /Tv  .z�@     �S  �O  /Us /Tv /Q0 0��@     �S  /Us /Tv /Q1  .c�@     �S  �O  /Uw /Ts  .��@     �S  	P  /U@/T6/Q0 .��@     �S  !P  /U~  .��@     �S  9P  /U}  .�@     �S  QP  /U}  ..�@     �S  iP  /U}  .j�@     �S  �P  /U}  .��@     �S  �P  /U}  .��@     �S  �P  /U}  .�@     �S  �P  /Us /Tv  .�@     �S  �P  /Us /Tv /Q0 0?�@     �S  /Us /Tv   5�k �3Q  6�v �rN  7res ��D   1c *�D  ��@     	      ��R  2>} +�/  �w �w 2L� ,�  'x x 2`5 -�  �x �x 2��  .�  z �y 2k /�   +{ { 2��  0�   �{ �{ 3�k 2�  g| ]| 3%k 3�  �| �| .��@     T  R  /Us /Tv  .��@     T  1R  /Us /Tv  .��@     T  OR  /Us /Tv  .4�@     T  mR  /Us /Tv  .K�@     T  �R  /Us /Tv  .j�@     T  �R  /Us /Tv  .|�@     T  �R  /Us /Tv  0��@     T  /Us /Tv   8Q  ��@     �       ��S  9Q  Y} O} :&Q  �} �} ;Q  P  hS  9Q  !~ ~ <P  =&Q  .�@     T  SS  /Us  >$�@     #T  /TC   .��@     3Q  S  /X0 0��@     #T  /TF  ?Vb Vb `?� � 6?3b 3b G?tk tk D?lk lk O?Nk Nk U	?l l T	?Ic Ic \	?�k �k X?�k �k I??k ?k �	?c c H?� �  6 �Y   �c  S#  �l �*  �@           �U Zs  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �  
K   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
K   /  ��   [r  �4 #�  �   �X  5�  
K   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K&  
�   P�  =_  ��   R�  N�  ��  ��   �p  W�  
K   3�  ��   ({  ��  ğ   F]  8�  
K   Y@  ��   �c  |  ��  l  ��  �   m c  
K   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {L  
K   ��  &�   �  º  GY  �f  ��   v�  ��  
K   �!  GQ   ϼ  �  �_  X  &�  �b   
K   �L  Cl [l 4�l h�l 4 �   W   	Y�  	%L  	��  	&L  ) 
{  J @
  � 
"�    � 
'
  �� 
*	�   
 
-  �9 
0	�    Ml  
3	�   $	
 
8	�   (C� 
;	�   ,� 
?	�   0� 
BR   8 �     =    o   
H	_  � 
K�    C� 
N	�   "8 
QR   t 
TR    . 
V!  k  }  R    r  	: 
��   	3 
��   	� 
��   	� 
��   	O 
��   	�
 
��   o  �   	R �  _  �   	� �  
K   r�  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	"|  *y  	��  +y  	I�  ,y  	�a  -y  B  �  =    4  �  =    
�	3	  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x ��   	�	  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4?	  �  �	   �	  �	  	��  My  	(h  N�   	l�  N�   	l
  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %
  l
  �
  =    	S�  'x
  t�   �   �
  �
  �
  =   �' �
  	��  1�
  	]  4�
  �
  �
  �
  =   � �
  	Zy  8�
  �    =   =   � �
  	��  ;  Ʃ  QK   "  .  D  =     3  	�  WD  �p  #�	  S�  $}  T}  %y    �  R   R    '	�  acv )U  ��  *a  ��  +m   �y -�  �Y  6�  ��  :
  s�  <
   �H  =
  xz  >�   �  x @�  
K   m  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �  
K   � )  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  uy  (x	z)   �u zm    � {	�    s |	�    � ~�   N�   )   ��  �	�    ��  �	�     J]  �)  z)  �)  =   � !�^  ��)  !�  �L  "K   ��,  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �)  \	X.   �Y  	�     *O  	�    ��  	�    �  	�    b�  	�    ��  	�    �  	�    +�  	�    Zp  	�     o�   	�   $ m�  !	�   ( 4�  "	�   , �  #	�   0 �  $	�   4 ��  %	�   8 L� &	�   < ��  '	�   @   (	�   D ��  )	�   H \q *	�   L z�  +	�   P �  ,	�   T /�  -	�   X ʤ  /-  X.  u.  =   � !��  1e.  
K   7�.  {�   U�  ~�   >	�.  �� @�.   s A
�   sx B�
  sy C�
   z)  Nz E�.  
K   p�/  �! 9& +! v( %# 0  B& @�! ��"  w#  	$  �-  S%  �)   0  @&  ��"    !0    m0    b-    �.    �$     /   @ %   � <"    U-    5'    	!  �]  ���1  `e �   x ��
  y ��
  z ��
   ��  ��1  (cN  ��1  0Mp �"  8�u �m  <� ��   @�H  ��1  Hr�  ��1  P��  ��1  X��  ��
  `m�  ��
  d��  ��
  h  ��
  l3F  ��
  p8F  ��
  t=F  ��
  x��  ��   |*� ��,  �y� ��1  �s ��   ��� ��.  ��  ��   ��  ��   �ʺ  ��   ��l  ��   �  �  �1  � ��  �   � ��  	�   � �R  �3  � f�  �   � I}  3	  � ��  �1  � �/  Gx  ��1  >} ��<   �}  �B  �|  �B  
 �1  X.  #d  HN�3  mo P)4   ��  Q�3  cmd R�	  �  W�
  (_  Y�
   #_  [�
  $bob ]�
  (�  a�   ,�[  b�   0sb  d�   4d]  g/4  8�W  h?4  P��  iy  h�� lO4  l�N  m�  |E�  p�  ��W  r_4  �~�  sO4  �*� tO4  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �)4  �$�R  ��    $��  ��   $�  ��   $h  �o4  $I�  �y  @ �1  �z �/  
K   1�3  ��   ��  ��   �y  9�3  
K   @)4  el �l �l  �3  �   ?4  =    y  O4  =    �   _4  =    y  o4  =    �.  4  =    hy ��1  (�	�4  in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
O4  �a  �
�   $ ��  ��4  ��	�5  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��5  ( �4  �5  =    ޴  ��4  	�  .y  	�  /y  	�  0y  	�  2y  	w�  8  	�  9�  	�  :�  	�_  ;�   	��  >y  	�  Jy  	"�  R�  	t�  S�   	�w  T�   	؜  Y�   	q�  [y  	Ƚ  ^�  	�  _�   	�y  `�   	b�  c�   	+�  fy  	��  iy  	֘ l�   	�J  x�   	��  y�   	ks  �   	�  ��   	J�  ��   	�i  ��   	��  �y  	��  �y  	��  �y  	<� �y  	��  �y  	��  �y  	5�  �y  	<m  ��   	 K  ��   	�R  ��   	op  ��   	�m  ��   	D  ��   	X�  ��   	If  ��   	� ��   	��  �y  	�U  �y  	`  �y  	J�  �y  	��  �y  	� ��  4  8  =    	�  �8  y  48  =    	� �$8  3	  P8  =   	 	,�  �@8  	R�  �h8  3	  3	  ~8  =    	�u  �n8  	��  ��5  	�e  ��   �   �8  =   � 	(�  ��8  	�  �y  !��  �  !�v  �   !n�  �   !4�  �   !*b �   !��  �	  H#	q9  � '
q9   �^  (1    .�  )	�   (o�  -1   0i�  .	�   8��  /
�9  < �   �9  =    �   �9  =    �  09  	��  .�9  	��  ��   	�\  �y  	�  ��9  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  ��	  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	�:  x E�
   y F�
   �{ Hd:  (T	�:  `e V   x W�
  y X�
  z Y�
    	�  [�:  �a	�;  = c�
   F�  d�
  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  o)4  ��  r
O4   iK  u�:  0��  x
�   XS�  {)4  `��  ~R   h��  ��   pu| �n<  x �}  X�n<  v1 �#=   v2 �#=  dx ��
  dy ��
  �  �B  �k �B  tag �B  �W  ��  �o �)=  $��  �=  4SX  ��<  8d�  ��<  @��  �
�   H��  �R   P t<  �;  �z ��:  �	�<  2�  ��
   ]  ��
  �h  �B  �N  �B  
�K  �B  >} ��<   z<  �}  ��<  
K   �=  ��   �  o�  ��   ��  ��<  �:  �
  9=  =    �u  ��;  �z ��1  8�	�=  v1 �#=   v2 �#=  82  ��
  Mp �"  [�  ��=   �  ��=   SX  ��<  (d�  ��<  0 �<  9=  A{ �Q=  4	2>  %x �
   %y 	�
  %dx 
�
  %dy �
   �o 2>   )�  �  0 �
  H>  =   =    (} �=  �  *�  &v  @2?   @�  4?   %x1 5�   %x2 6�    .]  8�
   5]  9�
   �� :�
   ��  =�    �  @�
    ��  C�
  $ �n  G?  ( 9x  H?  0 �^  I?  8 �=  B  >�  Kb>  &�h  PR@   s�  U@    �H  V@  %x1 X�   %x2 Y�   %gx \�
  %gy ]�
  %gz `�
   %gzt a�
  $ �x  d�
  ( � f�
  , ~�  i�
  0 t  k�
  4 .� l�   8 �  p@  @ 	�  r�   H 0?  U>  �h  t0?  �	Z@   �c  �y    �O  �Z@   �x  �
j@   B  j@  =    �  z@  =    I�  �%@  �	�@   �  ��     �  ��@   z@  �  ��@  '��	kA     ��
    �  �	�    t�  �	�    ��  �	�    /�  �	�    �  �	�  %top �	kA  (��  �	�  U(��  �	�  V(� �	kA  W(�  �	�  � �  |A  =   ? ��  ��@  	.L  &�A  �
  	׮  )�A  	�  +�A  	�  ,�A  	�Q  .@  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7B  �   	��  8B  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u FUB  �@  	��  H�   	��  I#=  	��  K�   	a� L?  	w�  N�   	P{ O�<  	��  Q�   	��  R�B  E=  	��  T�   	�� U�B  H>  	�}  W�   	u| X�=  	M�  Z�   	P�  [�=  	��  a�
  	��  b�
  	�  c�
  	�p  e"  	�T  fKC  4  	�a  j"  �   nC  =   � 	ը  l]C  "  �C  =   @ 	�p  mzC  	 �  p�
  	p|  q"  	$Y  v�   	�K  y�   	g  {�C  |A  	d�  |�C  	��   �
  		�  !�
  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�
  	`�  ,�
  	A�  -�
  	��  /�   	��  1�   	P�  2�   @  �D  =   =   / 	��  EuD  @  �D  =   / 	Ԁ  F�D  @  �D  =   =    	7� G�D  	�R  I�   	��  J@  	��  U�   	P�  \l  	��  ]l  	L�  ^l  	ߵ  _l  	�  al  	@�  ?  	[�  �=  	 �  �=  	SX  �<  	d�  �<  	��  �   	_�   �   	��  "y  	��  %y  	'�  &y  	�]  (y  #?  �E  =   � 	�P  *�E  	ӯ  +�E  #?  	|  -�E  @  	��  .�E  	��  /�E  F  'F  �   �    	��   ?  �    F  	qY   "3F  	�   #3F  B  hF  =   ? 	��   %WF  	��   &WF  �
  �F  =   � 	@Y   (�F  �
  �F  =   ? 	V�   )�F  @  �F  =    	�h  !�F  	�  !�F  @  	�  !@  	�f  !!WF  	r�  !"WF  	��  !%?  	��  !&?  	׆  !'�
  	��  !(�
  	�  !*�
  	��  !+�
  	�  "@  	��  "�   	�_  "�   	�_  "�   	b  "�
  	t  "�
  	j�  ""�	  	�  ":�   	��  ";�   	��  "<�   	�W  ">@  	hn  "@�
  	U~  "A�
  	�  "B�
  	 �  "C�
  	%�  "F�	  	�u  "H�	  	z  "I�	  	ʓ  #C  3	  GH  =    	��  #b7H  �   cH  =    	��  #cSH  	0K  #d�   	?�  #e�   #�	�H  x #��
   y #��
  dx #��
  dy #��
   ��  #��H  #��H  �p #�
)4  ��  #�
�=   #�	I  {q #��
   ��  #�y  d #�	�H   t�  #��H  I  8I  =   � 	r #�(I  	�T  #�PI  I  	l�  #��
  	�  #��
  	?k  #��
  	�d  #��
  	2~ #��H  	��  #�y  	��  #��
  	k�  #��
  	Z�  #��=  �=  �I  =    	�v  #��I  	�v  #��   	"�  #�)4  !�  #�	  !�U  #?  !��  #?  !t�  #�   !�  #	�   !.Y  #
�
  !7Y  #�
  !�h  #^J  )4  !*� #O4  !<i  #O4  	G  $y  	��  $�   
K   $��J  )top  �G  �  �]  $��J   $�	K  ��  $��=   ��  $��J  O{  $�
�   ��  $�
�   iK  $�K   �:  ��  $��J  K  0K  =    	��  $� K  "K   $cK  )up  �  �F  �S   FT  $
<K  "K   $�K  ��   �x  H�  ��  �H   ��  $pK  H$	^L   `e $    >} $�<   L� $�
   %low $�
  $ +� $ �
  ( �Z $!
�   , r� $"
�   0 �f  $#cK  4 �f  $$cK  8 ��  $%y  <%tag $&
�   @ *� $'�K  D �w $)�K  {L  {L  =    ^L  !�  $2kL  "K   $��L  ��   �s  z�  ��  �T  ܭ   gY  $��L  H$�	fM   `e $�    *� $��L   >} $��<    �W  $��
  ( �}  $��
  , L� $��
  0 ��  $�y  4 ��  $�
�   8%tag $�
�   < ��  $�
�   @  w $��L  �M  �M  =    fM  !j�  $sM  	 %V�   *dJ  2	�[e     *qJ  3	p[e     +dj -�@           �O  , �  )4  n~ Z~ ,	m )4  S E ,m�  )4  � � ,\q 	�   � ݀ -ang K   o� k� .�l 
�   �� �� .�R  KC  �� � .�l �
  G� C� .v� 
�   � }� /��@     Y  /�@     Y  09�@     $Y  �N  1U  0L�@     $Y  �N  1U  0:�@     0Y  $O  1U(1T:1Qv dv  $I"$,( 1$#( 2e�@     O  DO  1U�Q1T�U /j�@     Y  0��@     <Y  iO  1Us  3�@     <Y  1U�U  +am �x�@     �      �GP  ,m�  �)4  �� �� , �  �)4  �� � .�[ ��,  F� D� -mo �)4  k� i� /g�@     HY  /��@     TY  0��@     <Y  #P  1Us  /��@     Y  4!�@     `Y  1Q@K$  +7m M&�@     R      ��U  ,�k N)4  � �� ,m O)4  0� �� .�R  QKC  ь ό -i R
�   �� �� .� S�
  `� \� .*u T
�   ԍ �� 5V  q�@      �  m#Q  6:V  m� k� 7.V  8�  9FV  �� ��   5V  ��@        sdQ  6:V  �� �� 7.V  8  9FV  �� ސ   :�U  ��@      ��@            ��Q  6�U  � � 7�U   5�U  ��@      @  �R  6�U  -� +� 7�U  ;�U  P  6�U  S� Q� 7�U  4��@     SV  1Uu 1Td   :�U  ��@      ��@            �<R  6�U  y� w� 7�U   :�U  �@      �@            �vR  6�U  �� �� 7�U   :�U   �@       �@            �R  6�U  ő Ñ 7�U   :�U  >�@      >�@            �R  6�U  � � 7�U   0�@     V  S  1Uu 1Tt  0��@     �U   S  1Uu  0D�@     SV  =S  1Uu 1T: 0i�@     SV  ZS  1Uu 1TI 0t�@     hW  wS  1Us 1T0 0��@     hW  �S  1Us 1T01Q5 0��@     hW  �S  1Us 1T31Q1 0��@     hW  �S  1Us 1T31Q5 0�@     hW  �S  1Us 1T21Q1 0C�@     hW  !T  1Us 1T21Q5 0m�@     hW  CT  1Us 1T11Q1 0��@     hW  eT  1Us 1T11Q5 0��@     hW  �T  1Us 1Tv1Q1 0�@     �V  �T  1Us 1T61Q0 07�@     �V  �T  1Us 1T3 0^�@     �V  �T  1Us 1T71Q0 0��@     �V  U  1Us 1T41Q0 0��@     �V  -U  1Us 1T51Q0 0��@     �V  JU  1Us 1T2 0�@     �V  gU  1Us 1T8 0'�@     lY  �U  1U	P�B      0E�@     xY  �U  1U|  3r�@     �Y  1U0  <#m y  �U  =�R  KC  =�l �    +tl ��@            �V  >�R  KC  U>�|  
@  T ?�l �y  SV  @�R  �KC  @sb  ��   Aol �
�    B8l �y  Q�@     )       ��V  C�R  �KC  UDnum ��   � �  Bl �y  M�@           �hW  E�R  �KC  R� L� E~�  ��  �� �� Em �y  e� Y� F�l �y  � � FVm �y  � � 0��@     hW  6W  1Us  0��@     �Y  SW  1U01T! 4�@     hW  1Us   ?�l By  �W  @�R  CKC  @~�  D�  Gnum E�   A/m G
�    HhW  �@     1      �[X  6yW  X� P� 6�W  �� �� 6�W  *� � 9�W  �� �� IhW  �  9X  6�W  ӕ ѕ 6�W  �� �� 6yW  � � 8�  J�W    4B�@     lY  1U	��B     1Tv   HV  z�@            ��X  K.V  UK:V  T9FV  B� @�  H�U  ��@     x       �Y  K�U  U6�U  m� e� L�U  ��@            6�U  і ϖ 6�U  �� �� 4�@     SV  1Uu 1Td   MEf Ef xM� � &!Md  d  "	M�D �D '9M�e �e #s	MNl Nl #PM�b  �b  +M�( �( #kM��  ��  '7M11 11 #qM� � %6 mI   "h  S#  n �*  0�@     �      Pf �v  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  
K   "f  ��  WH  �~  �O  �m  ��   �  ��  ��  	 0t  r  e2    �0  }  ��  f  
K   J�  D   �C  
D  ���� �C  N�  ڵ  R�  �  
K   k,  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {�  
K   �k  &�   �  º  GY  �f  ��   v�  �8  t�  	 �   w  �  �  =   �' �  	��  
1�  	]  
4�  �  �  �  =   � �  	Zy  
8�  �  �  =   =   � �  	��  
;�  Ʃ  
QK       '  =       	�  
W'  �p  #D  J  Q   S�  $]  c  n  R    T}  %z  �  �  R   R    '	�  acv )8  ��  *Q  ��  +n   �y -�  �Y  6�  ��  :  s�  <   �H  =  xz  >�   �  x @�  �  -  =    y  =  =    
�	�  x ��   y ��  Mp ��  *� ��  ޽  ��   ~x �=  
K   �  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  
K   �t!  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�  (x	�!  �u z�   � {	�   s |	�   � ~�  N�  t!  ��  �	�   ��  �	�     J]  ��!  �!  "  =   � �^  ��!  �   $"   �  �"   K   �}%  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  1"  \	�&  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /�%  �&  �&  =   � ��  1�&  �]  ���(  `e �   x �w  y �w  z �w   ��  ��(  (cN  ��(  0Mp �  8�u ��  <� ��   @�H  ��(  Hr�  ��(  P��  �)  X��  �w  `m�  �w  d��  �w  h  �w  l3F  �w  p8F  �w  t=F  �w  x��  ��   |*� �}%  �y� �)  �s ��   ��� �)  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  �(  ���  �   ���  	�   ��R  �*  �f�  �   �I}  �  ���  �(  � '  Gx  �)  >} �b.   �}  ��  �|  ��  
 �(  �&  �!  !d  HN�*  mo P-   ��  Q�4  cmd Ra4  �  Ww  (_  Yw   #_  [w  $bob ]w  (�  a�   ,�[  b�   0sb  d�   4d]  g�4  8�W  h�4  P��  i�  h�� l"-  l�N  m,  |E�  p,  ��W  r�4  �~�  s"-  �*� t"-  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �-  �"�R  ��    "��  ��   "�  ��   "h  ��4  "I�  ��  @ $)  �z '  �  	��  ��   	�\  ��  	�  �;+  �  	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  �+  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	�+  x Ew   y Fw   �{ H�+  (T	6,  `e V   x Ww  y Xw  z Yw    	�  [�+  �a	-  = cw   F�  dw  �~ e�  h�  f�  
t�  g�  �k h�  tag i�  �N  l
�   ��  o-  ��  r
"-   iK  u6,  0��  x
�   XS�  {-  `��  ~R   h��  ��   pu| ��-  x +  �   2-  =    �}  X��-  v1 ��.   v2 ��.  dx �w  dy �w  �  ��  �k ��  tag ��  �W  �  �o ��.  $��  ��.  4SX  �b.  8d�  �b.  @��  �
�   H��  �R   P �-  2-  �z �B,  �	b.  2�  �w   ]  �w  �h  ��  �N  ��  
�K  ��  >} �b.   �-  �}  �
.  
K   ��.  ��   �  o�  ��   ��  �t.  �+  w  �.  =    �u  �2-  �z ��(  8�	E/  v1 ��.   v2 ��.  82  �w  Mp �  [�  �E/   �  �K/   SX  �b.  (d�  �b.  0 h.  �.  A{ ��.  4	�/  #x w   #y 	w  #dx 
w  #dy w  �o �/  )�  -  0 w  �/  =   =    (} ]/  �  *�  $v  @2�0  @�  4�0   #x1 5�   #x2 6�   .]  8w  5]  9w  �� :w  ��  =�   �  @w   ��  Cw  $�n  G�0  (9x  H�0  0�^  I�0  8 Q/  �  >�  K�/  $�h  PR�1  s�  U�1   �H  V�1  #x1 X�   #x2 Y�   #gx \w  #gy ]w  #gz `w   #gzt aw  $�x  dw  (� fw  ,~�  iw  0t  kw  4.� l�   8�  p�1  @	�  r�   H �0  �/  �h  t�0  �	�1  �c  ��   �O  ��1  �x  �
�1   �  �1  =    �  �1  =    I�  ��1  �	22  �  ��    �  �22   �1  �  �2  %��	�2    �w   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  #top �	�2  &��  �	�  U&��  �	�  V&� �	�2  W&�  �	�  � �   3  =   ? ��  �E2  	e3  ~�  k   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %3  e3  �3  =    	S�  'q3  >	�3  �� @)   s A
�   sx Bw  sy Cw   Nz E�3   	a4  ��  "�   E�  #�  e% $�  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�3  
K   1�4  ��   ��  ��   �y  9m4  �   �4  =    �  �4  =    �  �4  =    �3  �4  =    hy �$)  	.L  &�4  w  	׮  )�4  	�  +�4  	�  ,�4  	�Q  .�1  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7d5  �   	��  8d5  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�5  82  	��  H�   	��  I�.  	��  K�   	a� L�0  	w�  N�   	P{ Ob.  	��  Q�   	��  R6  �.  	��  T�   	�� U66  �/  	�}  W�   	u| XK/  	M�  Z�   	P�  [E/  	��  aw  	��  bw  	�  cw  	�p  e  	�T  f�6  �4  	�a  j  �   �6  =   � 	ը  l�6    �6  =   @ 	�p  m�6  	 �  pw  	p|  q  	$Y  v�   	�K  y�   	g  {07   3  	d�  |07  	��   w  		�  !w  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +w  	`�  ,w  	A�  -w  	��  /�   	��  1�   	P�  2�   �1  �7  =   =   / 	��  E�7  �1  8  =   / 	Ԁ  F�7  �1  &8  =   =    	7� G8  	�R  I�   	��  J�1  	��  U�   '	P�  \c8  V8  	��  ]c8  	L�  ^c8  	ߵ  _c8  	�  ac8  	@�  �0  	[�  E/  	 �  K/  	SX  b.  	d�  b.  	��  �   	_�   �   	��  "�  	��  %�  	'�  &�  	�]  (�  �0  -9  =   � 	�P  *9  	ӯ  +E9  �0  	|  -W9  �1  	��  .W9  	��  /W9  {9  �9  �   �    	��  �0  �   u9  	qY  "�9  	�  #�9  �  �9  =   ? 	��  %�9  	��  &�9  w  �9  =   � 	@Y  (�9  w  :  =   ? 	V�  ) :  �1  -:  =    	�h  :  	�  E:  �1  	�  �1  	�f  !�9  	r�  "�9  	��  %�0  	��  &�0  	׆  'w  	��  (w  	�  *w  	��  +w  	�  �1  	��  �   	�_  �   	�_  �   	b  w  	t  w  	j�  "+  	�  :�   	��  ;�   	��  <�   	�W  >�1  	hn  @w  	U~  Aw  	�  Bw  	 �  Cw  	%�  F+  	�u  H+  	z  I+  	ʓ  C  �  �;  =    	��  b�;  �   �;  =    	��  c�;  	0K  d�   	?�  e�   �	#<  x �w   y �w  dx �w  dy �w   ��  ��;  �Q<  �p �
-  ��  �
K/   �	�<  {q �w   ��  ��  d �	/<   t�  �Q<  �<  �<  =   � 	r ��<  	�T  ��<  �<  	l�  �w  	�  �w  	?k  �w  	�d  �w  	2~ �#<  	��  ��  	��  �w  	k�  �w  	Z�  �K/  K/  6=  =    	�v  �&=  	�v  ��   	"�  �-  �  +  �U  �0  ��  �0  t�  �   �  	�   .Y  
w  7Y  w  �h  �=  -  *� "-  <i  "-  	G  �  	��  �   0y	E>  `e {   >} |b.  r� }
�    �m ~
�   $�n 
�   ( �m ��=  8�	�>  `e �   >} �b.  r� �
�    �m �
�   $�n �
�   (�m �
�   ,�n �
�   0 qz �Q>  8�	'?  `e �   >} �b.  r� �
�    �n �
�   $�m �
�   (;n �
�   ,�n �
�   0 �w ��>  0�	~?  `e �   >} �b.  �n �
�    �m �
�   $��  �
�   ( �x �3?  
K   ��?  (top  �G  �  �]  ��?   �	@  ��  �K/   ��  ��?  O{  �
�   ��  �
�   iK  �@   6,  ��  ��?  @  $@  =    	��  �@   K   W@  (up  �  �F  �S   FT  
0@   K   �@  ��   �x  H�  ��  �H   ��  d@  H	RA  `e    >} b.  L� w   #low w  $+�  w  (�Z !
�   ,r� "
�   0�f  #W@  4�f  $W@  8��  %�  <#tag &
�   @*� '�@  D �w )�@  oA  oA  =    RA  �  2_A   K   ��A  ��   �s  z�  ��  �T  ܭ   gY  ��A  H�	ZB  `e �   *� ��A  >} �b.   �W  �w  (�}  �w  ,L� �w  0��  ��  4��  �
�   8#tag �
�   <��  �
�   @  w ��A  wB  wB  =    ZB  j�  gB  )Jn N�@     U       � C  *>} N$b.   � � +g P C  p� l� ,��@     (I  �B  -U0-T6-Q0 ,��@     4I  C  -Us  .��@     @I  -Uv   ~?  /!n 3@C  0g 3 C   )^n �@     p       �D  *��  	K/  �� �� *�m 
�   �� �� +i 
�   4� 2� +j 
�   [� W� 1>} b.  �� �� 1v� b.  �� �� 1~m K/  ߘ ݘ .V�@     LI  -Ts   2�n ���@     n       ��D  3��  �"K/  � 
� 4i ��   d� \� 4j ��   ř Ù 4min ��   � � 5>} �b.  � � 5�k �b.  4� 2� 5~m �K/  Y� W� .��@     LI  -Ts   2mn �a�@     @       �PE  3��  �$K/  �� �� 5�k �
�   � ֚ 4sec �b.  h� f� ,t�@     XI  6E  -Uv -Ts  .��@     PE  -T#-Q0  2�m ���@     �       �F  3>} �b.  �� �� 3�m ��   � ݛ 3�n ��   5� /� 5�x �F  �� �� ,��@     (I  �E  -U8-T6-Q0 ,�@     4I  �E  -Us  ,)�@     @I  F  -Uv  6H�@     dI   '?  7n �>F  8�x � F   2lm us�@     d       ��F  3>} u#b.  �� �� 5�x w�F  � � ,��@     (I  �F  -U8-T6-Q0 ,��@     4I  �F  -Us  ,��@     @I  �F  -Uv  6��@     dI   �>  7�n [G  8�x ["�F   2(n =�@     T       ��G  3>} =$b.  M� G� 5Dn ?�G  �� �� ,<�@     (I  lG  -U0-T6-Q0 ,G�@     4I  �G  -Us  .b�@     @I  -Uv   E>  7�m '�G  8Dn '$�G  9�m )	�    :$F  0�@     +       �H  ;1F  U<$F  5�@     %       =1F  ՝ ӝ   :&C  [�@     M       �QH  ;4C  U<&C  h�@             =4C  �� ��   :�G  ��@     :       ��H  =�G  %� � >�G  <�G  ��@     .       =�G  �� �� ?��@     .       @�G  ؞ ֞ 6��@     dI     :�F  ��@     =       �(I  =�F  � �� A�F  �  =�F  h� b� 6�@     dI  6�@     dI    B� � 6B3b 3b GB�m �m eB�m �m jBVb Vb `B� � ! �i   �k  S#  �o �*  ��@     a      �n �x  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  9�  t�   �   
(  K   `  �L  M M �L  0t  l  e2    �0  }  ��  `  K   J�  D   �C  
D  ���� �C  N�  ڵ  R�  
�  	 	a  ��  	"z   E�  	#z  e% 	$�  u  	%
�  �8 	&
�  ��  	)
�  /b  	-
�  ��  	.	�   a  	2
�  �T  	3
�   Mx 	4�  s  K   
�  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  
(t  K   
/�  ��   [r  �4 #�  �   �X  
5�  K   
:g  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  
K  �   
P�  =_  ��   R�  N�  ��  ��   �p  
Ws  K   3�  ��   ({  ��  ğ   F]  8�  K   Y  ��   �c  |  ��  l  ��  �   K   ko  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {  K   ��  &�   �  º  GY  �f  ��   v�  �{  K   ��  GQ   ϼ  �  �_  X  &�  �b   	�  �   	q    �   4  "  =   �' 
  	��  1"  	]  4?  4  4  V  =   � 
E  	Zy  8V  �  }  =   =   � 
g  	��  ;}  Ʃ  QK   
�  �  �  =     
�  	�  W�  �p  #�  �  �   S�  $�  �  �  R    T}  %  	    R   R    '	G  acv )�  ��  *�  ��  +�   �y -  �Y  6G  ��  :�  s�  <�   �H  =�  xz  >S   _  x @_  �  �  =    s  �  =    
�	  x ��   y ��  Mp ��  *� ��  ޽  ��   ~x ��  K   j
  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �  K   ��#  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  uv
  (x	w$  �u zj
   � {	�   s |	�   � ~G  N�  �#  ��  �	�   ��  �	�     J]  �
$  w$  �$  =   �  �^  ��$  �   �$  !  �  ��$  "K   �(  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �$  \	`)  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /(  `)  })  =   �  ��  1m)  K   pj*  �! 9& +! v( %# 0  B& @�! ��"  w#  	$  �-  S%  �)   0  @&  ��"    !0    m0    b-    �.    �$     /   @ %   � <"    U-    5'    	!  �]  ��@,  `e ��   x �(  y �(  z �(   ��  �@,  (cN  �@,  0Mp ��  8�u �j
  <� ��   @�H  �@,  Hr�  �@,  P��  �{,  X��  �(  `m�  �(  d��  �(  h  �(  l3F  �(  p8F  �(  t=F  �(  x��  ��   |*� �(  �y� ��,  �s ��   ��� ��,  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  @,  ���  �   ���  	�   ��R  g.  �f�  �   �I}    ���  @,  � j*  Gx  �{,  >} ��1   �}  ��  �|  ��  
 F,  `)  w$  #d  HNg.  mo P�0   ��  Q�7  cmd Ra  �  W(  (_  Y(   #_  [(  $bob ](  (�  a�   ,�[  b�   0sb  d�   4d]  g�7  8�W  h�7  P��  i�  h�� l�0  l�N  mo  |E�  po  ��W  r�7  �~�  s�0  �*� t�0  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��0  �$�R  ��    $��  ��   $�  ��   $h  ��7  $I�  ��  @ �,  �z j*  �  	��  ��   	�\  ��  	�  ��.  �  	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  �z.  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	[/  x E(   y F(   �{ H;/  (T	�/  `e V�   x W(  y X(  z Y(    	�  [g/  �a	�0  = c(   F�  d(  �~ e�  h�  f�  
t�  g�  �k h�  tag i�  �N  l
�   ��  o�0  ��  r
�0   iK  u�/  0��  x
�   XS�  {�0  `��  ~R   h��  ��   pu| �[1  x m.  �   �0  =    �}  X�[1  v1 �2   v2 �2  dx �(  dy �(  �  ��  �k ��  tag ��  �W  ��  �o �2  $��  �2  4SX  ��1  8d�  ��1  @��  �
�   H��  �R   P a1  �0  �z ��/  �	�1  2�  �(   ]  �(  �h  ��  �N  ��  
�K  ��  >} ��1   g1  �}  �s1  K   �2  ��   �  o�  ��   ��  ��1  [/  (  &2  =    �u  ��0  �z �F,  8�	�2  v1 �2   v2 �2  82  �(  Mp ��  [�  ��2   �  ��2   SX  ��1  (d�  ��1  0 �1  &2  A{ �>2  4	3  %x (   %y 	(  %dx 
(  %dy (  �o 3  )�  �  0 (  53  =   =    (} �2  �  *�  &v  @24  @�  44   %x1 5�   %x2 6�   .]  8(  5]  9(  �� :(  ��  =�   �  @(   ��  C(  $�n  G
4  (9x  H
4  0�^  I
4  8 �2  �  >�  KO3  &�h  PR�4  s�  U�4   �H  V�4  %x1 X�   %x2 Y�   %gx \(  %gy ](  %gz `(   %gzt a(  $�x  d(  (� f(  ,~�  i(  0t  k(  4.� l�   8�  p�4  @	�  r�   H 4  B3  �h  t4  �	G5  �c  ��   �O  �G5  �x  �
W5   �  W5  =    �  g5  =    I�  �5  �	�5  �  ��    �  ��5   g5  �  �t5  '��	X6    �(   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  %top �	X6  (��  �	�  U(��  �	�  V(� �	X6  W(�  �	�  � �  i6  =   ? ��  ��5  	�6  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %v6  �6  �6  =    	S�  '�6  K   77  {�   U�  ~�   >	S7  �� @�,   s A
�   sx B(  sy C(   Nz E7  K   1�7  ��   ��  ��   �y  9_7  �   �7  =    �  �7  =    �  �7  =    S7  �7  =    hy ��,  (�	<8  in ��   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�0  �a  �
�   $ ��  ��7  ��	�8  2�  �
�    I�  ��  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��8  ( <8  �8  =    ޴  �H8  	.L  &	9  (  	׮  )	9  	�  +	9  	�  ,	9  	�Q  .�4  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7{9  �   	��  8{9  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�9  �5  	��  H�   	��  I2  	��  K�   	a� L4  	w�  N�   	P{ O�1  	��  Q�   	��  R/:  22  	��  T�   	�� UM:  53  	�}  W�   	u| X�2  	M�  Z�   	P�  [�2  	��  a(  	��  b(  	�  c(  	�p  e�  	�T  f�:  �7  	�a  j�  �   �:  =   � 	ը  l�:  �  �:  =   @ 	�p  m�:  	 �  p(  	p|  q�  	$Y  v�   	�K  y�   	g  {G;  i6  	d�  |G;  	��   (  		�  !(  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +(  	`�  ,(  	A�  -(  	��  /�   	��  1�   	P�  2�   �4  �;  =   =   / 	��  E�;  �4  <  =   / 	Ԁ  F<  �4  =<  =   =    	7� G'<  	�R  I�   	��  J�4  	��  U�   	P�  \m  	��  ]m  	L�  ^m  	ߵ  _m  	�  am  	@�  4  	[�  �2  	 �  �2  	SX  �1  	d�  �1  	��  �   	_�   �   	��  "�  	��  %�  	'�  &�  	�]  (�  4  ==  =   � 	�P  *-=  	ӯ  +U=  4  	|  -g=  �4  	��  .g=  	��  /g=  �=  �=  �   �    	��  
4  �   �=  	qY  "�=  	�  #�=  �  �=  =   ? 	��  %�=  	��  &�=  (  >  =   � 	@Y  (�=  (  !>  =   ? 	V�  )>  5  =>  =    	�h  ->  	�  U>  5  	�  5  	�f  !�=  	r�  "�=  	��  %
4  	��  &
4  	׆  '(  	��  ((  	�  *(  	��  +(  	�  �4  	��  �   	�_  �   	�_  �   	b  (  	t  (  	j�  "z.  	�  :�   	��  ;�   	��  <�   	�W  >�4  	hn  @(  	U~  A(  	�  B(  	 �  C(  	%�  Fz.  	�u  Hz.  	z  Iz.  	ʓ  C�    �?  =    	��  b�?  �   �?  =    	��  c�?  	0K  d�   	?�  e�   �	3@  x �(   y �(  dx �(  dy �(   ��  ��?  �a@  �p �
�0  ��  �
�2   �	�@  {q �(   ��  ��  d �	?@   t�  �a@  �@  �@  =   � 	r ��@  	�T  ��@  �@  	l�  �(  	�  �(  	?k  �(  	�d  �(  	2~ �3@  	��  ��  	��  �(  	k�  �(  	Z�  ��2  �2  FA  =    	�v  �6A  	�v  ��   	"�  ��0   �  z.   �U  
4   ��  
4   t�  �    �  	�    .Y  
(   7Y  (   �h  �A  �0   *� �0   <i  �0  	G  �  	��  �   �   B  =    K   �;B  )top  �G  �  �]  �B   �	�B  ��  ��2   ��  �;B  O{  �
�   ��  �
�   iK  ��B   �/  ��  �GB  �B  �B  =    	��  ��B  "K   �B  )up  �  �F  �S   FT  
�B  "K   "C  ��   �x  H�  ��  �H   ��  �B  H	�C  `e �   >} �1  L� (   %low (  $+�  (  (�Z !
�   ,r� "
�   0�f  #�B  4�f  $�B  8��  %�  <%tag &
�   @*� '"C  D �w )/C  �C  �C  =    �C   �  2�C  "K   �FD  ��   �s  z�  ��  �T  ܭ   gY  �D  H�	�D  `e ��   *� �FD  >} ��1   �W  �(  (�}  �(  ,L� �(  0��  ��  4��  �
�   8%tag �
�   <��  �
�   @  w �SD  E  E  =    �D   j�  �D  ) &E  J @�E  � "�    � '

B  �� *	�   
 -�E  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 E   H	�E  � K�    C� N	�   "8 QR   t TR    . V�E  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   E  YF  ! 	R  NF  �E  pF  ! 	�  eF  K    rI  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	 !V�   a  	��  "M�  	(h  "N�   	l�  "N�   	�  #.�  	�  #/�  	�  #0�  	�  #2�  	w�  #8�  	�  #9�  	�  #:g  	�_  #;�   	��  #>�  	�  #J�  	"�  #R�  	t�  #S�   	�w  #T�   	؜  #Y�   	q�  #[�  	Ƚ  #^�  	�  #_�   	�y  #`�   	b�  #c�   	+�  #f�  	��  #i�  	֘ #l�   	�J  #x�   	��  #y�   	ks  #�   	�  #��   	J�  #��   	�i  #��   	��  #��  	��  #��  	��  #��  	<� #��  	��  #��  	��  #��  	5�  #��  	<m  #��   	 K  #��   	�R  #��   	op  #��   	�m  #��   	D  #��   	X�  #��   	If  #��   	� #��   	��  #��  	�U  #��  	`  #��  	J�  #��  	��  #��  	� #��  �7  �K  =    	�  #��K  �  �K  =    	� #��K    �K  =   	 	,�  #��K  	R�  #�L      #L  =    	�u  #�L  	��  #��8  	�e  #��   �   XL  =   � 	(�  #�GL  	�  #��   ��  #�   �v  #�    n�  #�    4�  #�    *b #�    ��  #+I  *�o ?
2  	pJf     *bp @
�0  	@Jf     *�p A�   	�Jf     +tmx B
(  	�If     +tmy C
(  	xIf     ,A  H
	�Jf     ,A  J
	�Jf     ,A  K
	TJf     *�o L
(  	�Jf     ,*A  P
	�Jf     ,FA  U
	�If     ,RA  V	`Jf     -q Q
(  	�Jf     -pq R
(  	�Jf     -�o T
�2  	�Jf     -�n U
�2  	`If     - o W
�0  	HJf     -�p Y
(  	�Jf     -q Z
(  	pIf     .^A  5
	�Jf     -�q 6
�0  	XJf     -Ap :
(  	�Jf     -Yq <�   	�Jf     -�n =
(  	PJf     -�p ?
(  	tIf      �o B(   �q C(  -�p t
�0  	�Jf     -�p �
�0  	�Jf     -�q �
�0  	hIf     -q ��   	�Jf     -�q 
�  	|If     -�o 
�  	�Jf     /�p o�O  0ld o$�2  1�o qK   	�e     20�  rK   34p v�     5?k X�  �A     L       �`P  6>} Y�1  �� �� 6)o Z�  
� � 7x \
�   E� C� 7y ]
�   p� h� 8$A     bh  9Us 9T|9Q	T
A       :(q 	�  �P  ;�p #�0  4mo �0   <.h �`A     �       ��Q  6�q ��0  Ҡ Π 6m�  ��0  � � 6\q ��   L� H� 7x �
�   �� �� 7y �
�   � � 7xl �
�   � � 7xh �
�   7� 5� 7yl �
�   \� Z� 7yh �
�   �� � =S� �(  �� �� 8�A     bh  9U~9Ts 9Q	 A       :�p �	�  �Q  ;�p �#�0  4dx �(  4dy �(  2S� �(   <�o �A     G       ��R  6�R  ��:  � � =Mp �
�   "�  � 7x1 �(  G� E� 7y1 �(  l� j� 4x2 �(  4y2 �(  >`A     nh  9X19Y	�A       :ro v	�  �R  0in v'�@  2<p x
�    <f V�A     z       ��S  ?t1 W�0  �� �� 6Mp X�  � �� 6#�  Y(  m� g� 6�  Z(  Ǥ �� 6\q [�   !� � 7x2 ](  w� u� 7y2 ^(  �� �� >A     nh  9X39Y	��@       5cg ,(  �A     �       �KT  ?t1 -�0  ť �� 6Mp .�  � � 6#�  /(  �� �� 7x2 1(  � � 7y2 2(  � 	� @A     zh  *T  9U�U 8�A     nh  9X39Y	H�@       5jp �	�  ��@     �      �pW  ?in �)�@  >� .� 7x �(  �� � 7y �(  j� b� 7z �(  � ը ={q �(  i� c� 7li ��2  �� �� 7th ��0  � � =�  �(  .� (� =S� �(  �� w� =�o �(  � � =�q �(  � � A�p ���@     @��@     �h  uU  9Ts  @��@     �h  �U  9U@>$ @ A     �h  �U  9Tv  @( A     �h  �U  9Tv  @8 A     �h  �U  9Uv  BE A     �h  @n A     �h  �U  9Us  B| A     �h  @� A     �h   V  9T|  @� A     �h  8V  9T|  @A     �h  PV  9T|  @6A     �h  tV  9U| ~ "9T}  " BeA     �h  @{A     �h  �V  9T}  @�A     �h  �V  9T}  @�A     �h  �V  9UD?$ @�A     �h  �V  9T}  @�A     �h  �V  9T}  @�A     �h  W  9U}  BA     �h  @&A     �h  =W  9U~ 9T  @9A     �h  [W  9U~ 9T  8YA     �h  9Us   5�n K�  H�@     e      ��X  ?in K�@  L� :� 7li M�2  � � 7th N�0  8� 2� =�  O(  �� �� =�o P(  Ĭ �� =�q Q(  "�  � =S� R(  M� E� @v�@     �h  ;X  9Us  B��@     �h  @��@     �h  `X  9Tv  @��@     �h  xX  9Tv  B<�@     �h  @R�@     �h  �X  9T}  8n�@     �h  9T}   <�q �A     �      ��Z  ?mo ��0  �� �� =�p �(  ?� =� =p �(  h� b� =0o �(  �� �� =7o �(  � � =�n �(  � � =�o �(  N� L� =�o ��   y� q� A>o �/A     A�p 4A     @EA     ?\  �Y  9Us  ClA     ?\  �Y  9U�U @�A     nh  �Y  9U| 9Tv 9X19Y	��@      @�A     nh  .Z  9U���9Tv 9X19Y	��@      @A     nh  ^Z  9U| 9T 9X19Y	��@      BiA     �h  ByA     �h  @�A     ?\  �Z  9Us  B�A     �h  B�A     �h  B�A     t[  8�A     ?\  9Us   5�q �	�  ��@     �       �t[  ?in �)�@  � � 7li ��2  9� 7� A9q ���@     @��@     �h  G[  9U	��B      @��@     �h  _[  9Qs  8�@     �h  9Us   DDo c�[  0ld c�2  2<p e�   2�p g�  2�q h�  2Hp i�  2�n k(  22p l(   5o -	�  �	A     X       �?\  6�p -$�0  b� \� =|p /�  �� �� 8
A     �\  9Us   :\i ��  �\  ;�p ��0  0x �(  0y �(  2�p �(  2�p �(  2<p �
�   29p �
�   4ld ��2   :�" ��  @]  ;�p ��0  0x �(  0y �(  4xl ��   4xh ��   4yl ��   4yh ��   4bx ��   4by ��   2p �/:   5So 	�  ��@     �      �^  6�p !�0  � � =�p (  �� �� 2�� �  =\q �   R� N� BU�@     �h  @�@     �h  �]  9U�h B��@     �h  B<�@     �h  @j�@     �h  ^  9U�h B��@     i   E�o �	�  3^  Fld � �2   G;i ��  �A     p      ��_  H�p ��0  �� �� Ix �(  �  � Iy �(  q� g� Jxl ��   � � Jxh ��   � � Jyl ��   6� 4� Jyh ��   [� Y� Jbx ��   �� ~� Jby ��   �� �� Kp �/:  �� �� @ A     i  4_  9U 9T��� @�A     bh  b_  9Us 9T���9Q	hA      @�A     $i  z_  9U~  8�A     0i  9U~   Eo a	�  �_  L�p a!�0  M�p c(   N�_  hA     |       �&`  O�_  � � P�_  Q�_  �  O�_  q� k� R�  S�_  �� �� 8�A     �h  9R
'    N^  �A     �      �a  O'^  �� �� T^  FA     M      ]a  O'^  b� ^� UyO  �A     �A     �       	Ha  O�O  �� �� V�A     �       S�O  ڶ ض T�O  �A     7       +a  S�O  � �� @A     <i  a  9U	ϱB     9T1 8"A     Hi  9T	�e       8�A     Ti  9T	رB        8}A     �h  9Us   81A     `i  9U	pJf     9Ts   N�R  �A     e       �.b  O�R  A� 7� S�R  �� �� T�R  �A            b  O�R  �� �� V�A            P�R  8�A     li  9TQ   B�A     �h  B�A     �h  B�A     xi   N�Q   A     �       ��b  O�Q  -� %� P�Q  P�Q  P�Q  Q�Q     O�Q  �� �� R   S�Q  � ޸ S�Q  � � S�Q  B� <� @bA     �i  �b  9Uv  8�A     �h  9Uv     N�\  A     �      �Xd  O�\  �� �� O�\  � � O�\  b� ^� P�\  P�\  P]  P]  P]  P&]  S2]  �� �� T�\  �A     �       ;d  O�\  º �� O�\  � � O�\  � � V�A     �       S�\  <� 8� S�\  x� r� S]  ǻ �� S]  � � S]  c� _� S&]  �� �� P2]  @A     bh  d  9Us 9T~ 9Q	��@      8|A     �i  9Us 9T~ 9Q	�A        8^A     i  9U�T9T�Q  N?\  �A     e      ��e  OQ\  ټ Ӽ O^\  +� %� Oi\  �� w� Pt\  P�\  P�\  P�\  P�\  T?\  �A     ,      �e  Oi\  � � O^\  �� �� OQ\  ˾ ɾ V�A     ,      St\  � � S�\  ,� (� S�\  h� b� S�\  �� �� S�\  � � @�A     $i  ]e  9Us  @	A     0i  ue  9Us  @�	A     �h  �e  9Qv  @�	A     �h  �e  9U| 9T} 9Qv  8�	A     �i  9Qs    8�A     �\  9Us 9Tv 9Q~   N`P  T
A     �       �g  OrP  +� %� PP  T`P  �
A     \       �f  OrP  {� w� V�
A     \       SP  �� �� @�
A     �h  �f  9Us 9T09Q09R: @�
A     �i  �f  9R& B A     �h  BA     �h  BA     �h  BA     �h    @_
A     �[  �f  9Us  @}
A     �h  g  9Us 9T
 8�
A     �i  9Us   Nt[  ,A     �       �bh  O�[  �� �� P�[  P�[  P�[  P�[  P�[  P�[  Qt[  0  O�[  D� @� R0  S�[  �� }� S�[  �� �� S�[  �� �� S�[  � � S�[  R� P� S�[  y� u� @iA     �h  �g  9Qs  @{A     �i  �g  9U09T0 @�A     �i  h  9U09T0 B�A     �i  B�A     �h  @�A     �h  Kh  9U|  8 A     �h  9U|     W�h �h �	WSp Sp �W�e �e r	W�o �o 7WH_  H_  #	Wd  d  "	W�g �g �W�e �e vWcq cq wXdj dj W��  ��  $7W�q �q �W� � %!W�e �e s	X7m 7m W3, 3, �Wi i �W�d �d �W��  ��  %WSJ SJ &"	WF�  F�  bWbo bo �W� � !6W�i �i 1W�f �f �	WDq Dq �	W�q �q <W�( �( kW11 11 qWEf Ef xW�h �h �	 �X   �p  S#  �r �*  5A     `
      o� �|  �)  �=   ,	  int ^&  9�  t�   D   [   �   �   �L  M M �L  �  	�1  @  
Q     
�   	1   
62  #	1   
  &	1   
�5  )	1    
�@  ,	1   (
.  -	1   0
*  2D   8
;:  5D   < #  1  �K 8"�   �  KB  *  �  LB  �  MB  0t  l  e2    �0  }  ��  `  �   J�  D   �C  
D  ���� �C  N�  ڵ  R�  �  �   	   7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  	(�  �   	/Y  ��   [r  �4 #�  �   �X  	5,  �   	:�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  	Ke  D   	P  =_  ��   R�  N�  ��  ��   �p  	W�  �   
3:  ��   ({  ��  ğ   F]  
8  �   
Y  ��   �c  |  ��  l  ��  �   �   
k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  
{  �   
�  &�   �  º  GY  �f  ��   v�  
��  �   
�T  GQ   ϼ  �  �_  X  &�  �b   �  d  =    s  t  =    
�	�  x ��   y ��  
Mp ��  
*� ��  
޽  ��   ~x �t   	S  
��  "z   
E�  #z  
e% $�  
u  %
�  
�8 &
�  
��  )
�  
/b  -
�  
��  .	D   
a  2
�  
�T  3
�   Mx 4�  �  l   e  S  ��  M�  (h  ND   l�  ND   	�  
~�     
�S  
D   
��   
D   
  !
D   
�g  "
D   
�^  #
D    ��  %�  �    =    S�  '   g   -  =   �'   ��  1-  ]  4J  g   g   a  =   � P  Zy  8a  �  �  =   =   � r  ��  ;�  Ʃ  Q�   �  �  �  =     �  �  W�  �p  #l  S�  $�  �  �  K    T}  %      K   K    '	E  acv )�  ��  *�  ��  +�   �y -  �Y  6E  	��  :�  
s�  <�   
�H  =�  
xz  >Q   ]  x @]  �   �
  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  �   ��$  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u  (x	%  �u z�
   � {	D   s |	D   � ~E  N�  �$  ��  �	D   ��  �	D     J]  ��$  %   %  =   � �^  �%    8%    �  �-%  !�   ��(  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  E%  \	�)  �Y  	D    *O  	D   ��  	D   �  	D   b�  	D   ��  	D   �  	D   +�  	D   Zp  	D    o�   	D   $m�  !	D   (4�  "	D   ,�  #	D   0�  $	D   4��  %	D   8L� &	D   <��  '	D   @  (	D   D��  )	D   H\q *	D   Lz�  +	D   P�  ,	D   T/�  -	D   X ʤ  /�(  �)  *  =   � ��  1�)  �   76*  {�   U�  ~�   >	r*  
�� @r*   
s A
D   sx B[   sy C[    %  Nz E6*  �   pd+  �! 9& +! v( %# 0  B& @�! ��"  w#  	$  �-  S%  �)   0  @&  ��"    !0    m0    b-    �.    �$     /   @ %   � <"    U-    5'    	!  	�]  ��:-  
`e ��   x �[   y �[   z �[    
��  �:-  (
cN  �:-  0
Mp ��  8
�u ��
  <
� �D   @
�H  �:-  H
r�  �:-  P
��  �u-  X
��  �[   `
m�  �[   d
��  �[   h
  �[   l
3F  �[   p
8F  �[   t
=F  �[   x
��  �D   |
*� ��(  �
y� �{-  �
s �D   �
�� �r*  �
�  �D   �
�  �D   �
ʺ  �D   �
�l  �D   � �  :-  ���  D   ���  	D   ��R  [/  �f�  D   �I}  �  ���  :-  � d+  	Gx  �u-  
>} ��7   
�}  ��  
�|  ��  
 @-  �)  "d  HN[/  mo P�/   
��  Q�/  cmd RS  
�  W[   
(_  Y[    
#_  [[   $bob ][   (
�  aD   ,
�[  bD   0
sb  dD   4
d]  g�/  8
�W  h�/  P
��  i�  h
�� l�/  l
�N  m�  |
E�  p�  �
�W  r�/  �
~�  s�/  �
*� t�/  �
�� wD   �
��  xD   �
X�  |D   �
�e  D   �
��  �D   �
g  �D   �
�u  �D   �
|G �  �
Q  �D   �
�  �D   �
o�  ��/  �#�R  �D    #��  �D   #�  �D   #h  ��/  #I�  ��  @ �-  �z d+  �   1�/  ��   ��  ��   �y  9n/  a/  D   �/  =    �  �/  =    D   �/  =    �  �/  =    x*  �/  =    hy ��-  (�	a0  in ��   
d  �
D   
�x  �
D   
D  �
D   
5O  �
D   
�� �
�/  
�a  �
D   $ ��  ��/  ��	1  
2�  �
D    
I�  ��  
r�  �
D   
�H  �
D   
*F  �
D   
��  �
D   
	�  �
D   
ѵ  �
D   
��  �
D    
F� �
D   $
�  �1  ( a0  1  =    ޴  �m0  �  .�  �  /�  �  0�  �  2�  w�  8Y  �  9   �  :�  �_  ;  ��  >�  �  J�  "�  R  t�  SD   �w  TD   ؜  YD   q�  [�  Ƚ  ^  �  _D   �y  `D   b�  cD   +�  f�  ��  i�  ֘ lD   �J  xD   ��  yD   ks  D   �  �D   J�  �D   �i  �D   ��  ��  ��  ��  ��  ��  <� ��  ��  ��  ��  ��  5�  ��  <m  �D    K  �D   �R  �D   op  �D   �m  �D   D  �D   X�  �D   If  �D   � �D   ��  ��  �U  ��  `  ��  J�  ��  ��  ��  � �:  �/  �3  =    �  �z3  �  �3  =    � ��3  �  �3  =   	 ,�  ��3  R�  ��3  �  �  �3  =    �u  ��3  ��  �1  �e  �  #  %4  =   � (�  �4  �  ��  ��  :  �v  D   n�  D   4�  D   *b D   ��  r  ��  �  �\  ��  �  ��4  �  ��  �D   ��  �D   2�  ��  ��  �D   Ɇ  �_  ��  �D   ��  �D   �h  �D   rK  �D   l�  �D   ]�  �D   ��  �D   C	f5  x E[    y F[    �{ HF5  (T	�5  
`e V�   x W[   y X[   z Y[     	�  [r5  �a	�6  
= c[    
F�  d[   
�~ e�  
h�  f�  

t�  g�  
�k h�  tag i�  
�N  l
D   
��  o�/  
��  r
�/   
iK  u�5  0
��  x
D   X
S�  {�/  `
��  ~K   h
��  �D   p
u| �P7  x 	�}  X�P7  v1 �8   v2 �8  dx �[   dy �[   
�  ��  
�k ��  tag ��  
�W  �T  
�o �8  $
��  ��7  4
SX  ��7  8
d�  ��7  @
��  �
D   H
��  �K   P V7  �6  �z ��5  �	�7  
2�  �[    
]  �[   
�h  ��  
�N  ��  

�K  ��  
>} ��7   \7  �}  �h7  �   ��7  ��   �  o�  ��   ��  ��7  f5  [   8  =    �u  ��6  �z �@-  8�	�8  v1 �8   v2 �8  
82  �[   
Mp ��  
[�  ��8  
 �  ��8   
SX  ��7  (
d�  ��7  0 �7  8  A{ �38  4	9  $x [    $y 	[   $dx 
[   $dy [   �o 9  )�  d  0 [   *9  =   =    (} �8  �  *�  %v  @2�9  @�  4�9   $x1 5D   $x2 6D   .]  8[   5]  9[   �� :[   ��  =D   �  @[    ��  C[   $�n  G�9  (9x  H�9  0�^  I�9  8 �8  �  >�  KD9  %�h  PR�:  s�  U�:   �H  V�:  $x1 XD   $x2 YD   $gx \[   $gy ][   $gz `[    $gzt a[   $�x  d[   (� f[   ,~�  i[   0t  k[   4.� lD   8�  p�:  @	�  rD   H :  79  �h  t:  �	<;  �c  ��   �O  �<;  �x  �
L;   �  L;  =    �  \;  =    I�  �;  �	�;  �  �D    �  ��;   \;  �  �i;  &��	M<    �[    �  �	D   t�  �	D   ��  �	D   /�  �	D   �  �	�  $top �	M<  '��  �	�  U'��  �	�  V'� �	M<  W'�  �	�  � �  ^<  =   ? ��  ��;  .L  &w<  [   ׮  )w<  �  +w<  �  ,w<  �Q  .�:  ��  0D   ��  1D   (_  2D   դ  4D   �j  7�<  D   ��  8�<  @�  <D   �O  =D   (g  >D   �^  ED   �u F7=  �;  ��  HD   ��  I8  ��  KD   a� L�9  w�  ND   P{ O�7  ��  QD   ��  R�=  '8  ��  TD   �� U�=  *9  �}  WD   u| X�8  M�  ZD   P�  [�8  ��  a[   ��  b[   �  c[   �p  e�  �T  f->  �/  �a  j�  D   P>  =   � ը  l?>  �  m>  =   @ �p  m\>   �  p[   p|  q�  $Y  vD   �K  yD   g  {�>  ^<  d�  |�>  ��   [   	�  ![   �3 #D   _  $D   -�  (D   �f  )D   �G  +[   `�  ,[   A�  -[   ��  /D   ��  1D   P�  2D   �:  m?  =   =   / ��  EW?  �:  �?  =   / Ԁ  Fy?  �:  �?  =   =    7� G�?  �R  ID   ��  J�:  ��  UD   (P�  \�?  �?  ��  ]�?  L�  ^�?  ߵ  _�?  �  a�?  @�  �9  [�  �8   �  �8  SX  �7  d�  �7  ��  D   _�   D   ��  "�  ��  %�  '�  &�  �]  (�  :  �@  =   � �P  *�@  ӯ  +�@  :  |  -�@  �:  ��  .�@  ��  /�@   A  A  D   D    ��  �9  �   �@  qY  "A  �  #A  �  QA  =   ? ��  %@A  ��  &@A  [   yA  =   � @Y  (iA  [   �A  =   ? V�  )�A  �:  �A  =    �h  �A  �  �A  �:  �  �:  �f  !@A  r�  "@A  ��  %�9  ��  &�9  ׆  '[   ��  ([   �  *[   ��  +[   �  �:  ��  D   �_  D   �_  D   b  [   t  [   j�  "_  �  :D   ��  ;D   ��  <D   �W  >�:  hn  @[   U~  A[   �  B[    �  C[   %�  F_  �u  H_  z  I_  ʓ  C�  �  0C  =    ��  b C  D   LC  =    ��  c<C  0K  dD   ?�  eD   �	�C  x �[    y �[   dx �[   dy �[    ��  �pC  ��C  �p �
�/  ��  �
�8   �	D  
{q �[    
��  ��  d �	�C   t�  ��C  D  !D  =   � r �D  �T  �9D  D  %r �KD  QD  )�  `D  9D   l�  �[   �  �[   ?k  �[   �d  �[   2~ ��C  ��  ��  ��  �[   k�  �[   Z�  ��8  �8  �D  =    �v  ��D  �v  �D   "�  ��/  �  _  �U  �9  ��  �9  t�  D   �  	D   .Y  
[   7Y  [   �h  hE  �/  *� �/  <i  �/  G  �  ��  D   �   ��E  *top  �G  �  �]  ��E   �	F  
��  ��8   
��  ��E  
O{  �
D   
��  �
D   
iK  �F   �5  ��  ��E  F  :F  =    ��  �*F  !�   mF  *up  �  �F  �S   FT  
FF  !�   �F  ��   �x  H�  ��  �H   ��  zF  H	hG  `e �   >} �7  L� [    $low [   $+�  [   (�Z !
D   ,r� "
D   0�f  #mF  4�f  $mF  8��  %�  <$tag &
D   @*� '�F  D �w )�F  �G  �G  =    hG  �  2uG  !�   ��G  ��   �s  z�  ��  �T  ܭ   gY  ��G  H�	pH  `e ��   *� ��G  >} ��7   �W  �[   (�}  �[   ,L� �[   0��  ��  4��  �
D   8$tag �
D   <��  �
D   @  w ��G  �H  �H  =    pH  j�  }H  +`D  !		�Jf     +lD  "		�Jf     +xD  #		�Jf     +�D  $		�Vf     +!D  	 Kf     +-D  	�Jf     +�D  	�Vf     ,gr 
�  	�Jf     ,pr  D   	�Jf      s �[   �	�I  $len �	D    0�  �K   s ��   as �`I  �I  �I  =    -�r ��I  	@�B     .Sp ]�  3A     b      ��L  /x1 ^[   �� �� /y1 _[   � � /x2 `[   x� r� /y2 a[   �� �� 0�  b	D   � � 0�r cKD  V� R� 1xt1 e[   �� �� 1yt1 f[   $� "� 1xt2 g[   S� G� 1yt2 h[   �� �� 2�  j[   w� o� 2�  k[   �� �� 2Gr m[   2� $� 2xr o[   �� �� 2�r p[   � � 2r r
D   ?� ;� 2 r s
D   }� y� 2�r u
D   �� �� 2Rs v
D   � � 2r� x
D   x� n� 3A     �X  �K  4Us 4T~ O&~ '~ O& 3;A     �X  �K  4Us 4T~ O&~ '~ O& 3nA     �X  �K  4U 4T��� 5�A     �X  5�A     �X  3�A     �X  /L  4Ts  3A     &R  ]L  4U���4T} 4Q	OA      3"A     �Q  �L  4U���4T} 4Q	YA      6�A     {M  4U��4T@<$  7�r ;�L  8�q ;#D   8yr ;@9D  9;Q =	D    :Or 5A     t       �{M  0;Q )D   � �� 0�| 7D   i� c� 1i 	D   �� �� 282  D   $� � 2�8 	D   �� �� 20�  K   �  �  .�r ��  �A     s       �,N  0ڈ �?D  +� %� 0�r �[   }� w� 2r� �D   �� �� 2S� �[   I� G� 2s �9D  n� l� 1in �9D  �� �� ;A     4U|   .�r f	�  YA     �       ��O  0�p f)�/  �� �� 1x1 h[   5� 3� 1y1 i[   Z� X� 1x2 j[   � }� 1y2 k[   �� �� 1s1 mD   �� �� 1s2 nD   � � 2vs p�  *� (� <dl r�C  ��2{q t[   n� l� =�L  A     A            �{O  >�L  �� �� >�L  �� �� ?A            @�L  5A     DW    3�A     U  �O  4U~ 4T| 4Q	�Vf      3�A     U  �O  4U���4Ts 4Q	�Vf      A�A     T  4U	�Vf     4T��  .1r /�  OA     
      ��Q  /ld / �8  �� �� 1s1 1D   5� -� 1s2 2D   �� �� 2{q 3[   �� �� <dl 4�C  �P=�L  6A     6A            [�P  >�L  �� �� >�L  � � ?6A            @�L  5CA     DW    3�A     U  �P  4Q	�Vf      3�A     U  Q  4Q	�Vf      3�A     �V  5Q  4Qs  3�A     �V  MQ  4Qs  3�A     �T  kQ  4Uu 4Tt  A�A     T  4U	�Vf     4Tw   .�h ��  iA     W       �R  /x �	D   @� :� /y �	D   �� �� 0ڈ � R  �� �� 2y �/  G� E� ;�A     4Us   )�   R  �/   R  BDq ��  �A     }       ��R  /x �	D   p� j� /y �	D   �� �� 0ڈ ��R  � � 982  �D   2*  ��9  w� u� 1ld ��8  �� ��  )�  �R  �8   �R  C�d �4A     �       �rS  0�p ��/  �� �� 1ss ��=  ,� &� 1sec ��7  }� {� 2r �D   �� �� 9r �D   2
 �hE  
� � 5CA     �X   Ci V�A     �       ��S  D�p V$�/  U2r X
D   3� -� 9r Y
D    C�g ':A     Y       �T  D �  '�8  U2g� )�7  �� �� 2� *�7  �� ��  Es �[   �A     s       ��T  Fv2 ��T  � �� Fv1 ��T  �� v� G{q �[   VHnum �[   �� �� Hden �[   <� 4� 5�A     �X  5	A     �X  5A     �X  53A     �X  IEA     �X   �C  JDs ��A            �U  Kli ��8  UKdl ��T  T E/s �D   8A     �       ��U  Fx �[   �� �� Fy �[   �� �� L��  ��T  I� A� Hdx �[   �� �� Hdy �[   �� �� MϷ  �[   � � M�T  �[   C� A� 5�A     �X  A�A     �X  4Uv 8&  Ebo iD   jA     �       ��V  L[s jw<  l� f� Fld k�8  �� �� Hp1 m
D   P� 4� Hp2 n
D   �� �� 3A     �V  nV  4Q|  3A     �V  �V  4Q|  A,A     �V  4Q|   N�q =D   �V  Ox >[   Oy ?[   P��  @�8  Qdx B[   Qdy C[   RϷ  D[   R�T  E[    E�h ,[   �A     #       �DW  Fdx -[   6� ,� Fdy .[   �� ��  S�L  �A     1       ��W  >�L  3� -� >�L  �� �� T�L  �� �� 3�A     �L  �W  4Uy  3�A     �L  �W  4Uy 6�A     �L  4Uy  S�V  �A     m       ��X  >�V  �� �� >�V  9� 3� >�V  �� �� @�V  T�V  �� �� T�V  *� &� T�V  b� `� U�V  
A            �X  >�V  �� �� >�V  �� �� >�V  �� �� ?
A            @�V  @�V  @�V  @�V    5MA     �X  A[A     �X  4Uv   VH_  H_  #	Vd  d  "	V3, 3, � �^   v  S#  �s �*  �A     B      �� �  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �   	"  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�  4  
K   "z  ��  WH  �~  �O  �m  ��   �  ��  ��  	 
K   	�  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  	(z  
K   	/�  ��   [r  �4 #�  �   �X  	5�  
K   	:m  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  	K
  
�   	P�  =_  ��   R�  N�  ��  ��   �p  	Wy  
K   
3�  ��   ({  ��  ğ   F]  
8�  
K   
Y$  ��   �c  |  ��  l  ��  �   
K   
ku  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  
{$  
K   
��  &�   �  º  GY  �f  ��   v�  
��  
K   
��  GQ   ϼ  �  �_  X  &�  �b   t�   �   �      =   �' 
  	��  1  	]  48      O  =   � >  	Zy  8O  �  v  =   =   � `  	��  ;v  Ʃ  QK   �  �  �  =     �  	�  W�  �p  #�  �  �   S�  $�  �  �  R    T}  %�      R   R    '	@  acv )�  ��  *�  ��  +�   �y -  �Y  6@  ��  :�  s�  <�   �H  =�  xz  >L   X  x @X  B  �  =    4  �  =    
�	  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x ��  
K   c
  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �  
K   ��#  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  uo
  (x	p$  �u zc
   � {	�   s |	�   � ~@  N�  �#  ��  �	�   ��  �	�     J]  �$  p$  �$  =   �  �^  �}$  �   �$  !  �  ��$  "K   ��'  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �$  \	Y)  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /(  Y)  v)  =   �  ��  1f)  
K   pc*  �! 9& +! v( %# 0  B& @�! ��"  w#  	$  �-  S%  �)   0  @&  ��"    !0    m0    b-    �.    �$     /   @ %   � <"    U-    5'    	!  �]  ��9,  `e ��   x ��  y ��  z ��   ��  �9,  (cN  �9,  0Mp ��  8�u �c
  <� ��   @�H  �9,  Hr�  �9,  P��  �t,  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� ��'  �y� �z,  �s ��   ��� ��,  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  9,  ���  �   ���  	�   ��R  `.  �f�  �   �I}    ���  9,  � c*  Gx  �t,  >} ��1   �}  �B  �|  �B  
 ?,  Y)  p$  #d  HN`.  mo P~0   ��  Qy7  cmd R"  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g�7  8�W  h�7  P��  iy  h�� l�0  l�N  mu  |E�  pu  ��W  r�7  �~�  s�0  �*� t�0  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �~0  �$�R  ��    $��  ��   $�  ��   $h  ��7  $I�  �y  @ �,  �z c*  �  	��  ��   	�\  �y  	�  ��.  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  �s.  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	T/  x E�   y F�   �{ H4/  (T	�/  `e V�   x W�  y X�  z Y�    	�  [`/  �a	~0  = c�   F�  d�  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  o~0  ��  r
�0   iK  u�/  0��  x
�   XS�  {~0  `��  ~R   h��  ��   pu| �T1  x f.  �   �0  =    �}  X�T1  v1 �	2   v2 �	2  dx ��  dy ��  �  �B  �k �B  tag �B  �W  ��  �o �2  $��  ��1  4SX  ��1  8d�  ��1  @��  �
�   H��  �R   P Z1  �0  �z ��/  �	�1  2�  ��   ]  ��  �h  �B  �N  �B  
�K  �B  >} ��1   `1  �}  �l1  
K   ��1  ��   �  o�  ��   ��  ��1  T/  �  2  =    �u  ��0  �z �?,  8�	�2  v1 �	2   v2 �	2  82  ��  Mp ��  [�  ��2   �  ��2   SX  ��1  (d�  ��1  0 �1  2  A{ �72  4	3  %x �   %y 	�  %dx 
�  %dy �  �o 3  )�  �  0 �  .3  =   =    (} �2  �  *�  &v  @2�3  @�  4�3   %x1 5�   %x2 6�   .]  8�  5]  9�  �� :�  ��  =�   �  @�   ��  C�  $�n  G4  (9x  H4  0�^  I4  8 �2  B  >�  KH3  &�h  PR�4  s�  U�4   �H  V�4  %x1 X�   %x2 Y�   %gx \�  %gy ]�  %gz `�   %gzt a�  $�x  d�  (� f�  ,~�  i�  0t  k�  4.� l�   8�  p�4  @	�  r�   H 4  ;3  �h  t4  �	@5  �c  �y   �O  �@5  �x  �
P5   B  P5  =    �  `5  =    I�  �5  �	�5  �  ��    �  ��5   `5  �  �m5  '��	Q6    ��   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  %top �	Q6  (��  �	�  U(��  �	�  V(� �	Q6  W(�  �	�  � �  b6  =   ? ��  ��5  	�6  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %o6  �6  �6  =    	S�  '�6  
K   77  {�   U�  ~�   >	L7  �� @�,   s A
�   sx B�  sy C�   Nz E7  
K   1y7  ��   ��  ��   �y  9X7  
K   @�7  el �l �l  �   �7  =    y  �7  =    y  �7  =    L7  �7  =    hy ��,  (�	V8  in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�0  �a  �
�   $ ��  ��7  ��	�8  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��8  ( V8  9  =    ޴  �b8  	.L  &#9  �  	׮  )#9  	�  +#9  	�  ,#9  	�Q  .�4  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�9  �   	��  8�9  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�9  �5  	��  H�   	��  I	2  	��  K�   	a� L�3  	w�  N�   	P{ O�1  	��  Q�   	��  RI:  +2  	��  T�   	�� Ug:  .3  	�}  W�   	u| X�2  	M�  Z�   	P�  [�2  	��  a�  	��  b�  	�  c�  	�p  e�  	�T  f�:  �7  	�a  j�  �   �:  =   � 	ը  l�:  �  ;  =   @ 	�p  m;  	 �  p�  	p|  q�  	$Y  v�   	�K  y�   	g  {a;  b6  	d�  |a;  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   �4  <  =   =   / 	��  E<  �4  5<  =   / 	Ԁ  F%<  �4  W<  =   =    	7� GA<  	�R  I�   	��  J�4  	��  U�   	P�  \.  	��  ].  	L�  ^.  	ߵ  _.  	�  a.  	@�  �3  	[�  �2  	 �  �2  	SX  �1  	d�  �1  	��  �   	_�   �   	��  "y  	��  %y  	'�  &y  	�]  (y  	4  W=  =   � 	�P  *G=  	ӯ  +o=  	4  	|  -�=  �4  	��  .�=  	��  /�=  �=  �=  �   �    	��  4  �   �=  	qY  "�=  	�  #�=  B  �=  =   ? 	��  %�=  	��  &�=  �  >  =   � 	@Y  (>  �  ;>  =   ? 	V�  )*>  �4  W>  =    	�h  G>  	�  o>  �4  	�  �4  	�f  !�=  	r�  "�=  	��  %4  	��  &4  	׆  '�  	��  (�  	�  *�  	��  +�  	�  �4  	��  �   	�_  �   	�_  �   	b  �  	t  �  	j�  "s.  	�  :�   	��  ;�   	��  <�   	�W  >�4  	hn  @�  	U~  A�  	�  B�  	 �  C�  	%�  Fs.  	�u  Hs.  	z  Is.  	ʓ  C�    �?  =    	��  b�?  �   �?  =    	��  c�?  	0K  d�   	?�  e�   �	M@  x ��   y ��  dx ��  dy ��   ��  �@  �{@  �p �
~0  ��  �
�2   �	�@  {q ��   ��  �y  d �	Y@   t�  �{@  �@  �@  =   � 	r ��@  	�T  ��@  �@  	l�  ��  	�  ��  	?k  ��  	�d  ��  	2~ �M@  	��  �y  	��  ��  	k�  ��  	Z�  ��2  �2  `A  =    	�v  �PA  	�v  ��   	"�  �~0   �  s.   �U  4   ��  4   t�  �    �  	�    .Y  
�   7Y  �   �h  �A  ~0   *� �0   <i  �0  	G  y  	��  �   �   4B  =    
K   �UB  )top  �G  �  �]  �4B   �	�B  ��  ��2   ��  �UB  O{  �
�   ��  �
�   iK  ��B   �/  ��  �aB  �B  �B  =    	��  ��B  "K   C  )up  �  �F  �S   FT  
�B  "K   <C  ��   �x  H�  ��  �H   ��  C  H	�C  `e �   >} �1  L� �   %low �  $+�  �  (�Z !
�   ,r� "
�   0�f  #C  4�f  $C  8��  %y  <%tag &
�   @*� '<C  D �w )IC  D  D  =    �C   �  2	D  "K   �`D  ��   �s  z�  ��  �T  ܭ   gY  �,D  H�	E  `e ��   *� �`D  >} ��1   �W  ��  (�}  ��  ,L� ��  0��  �y  4��  �
�   8%tag �
�   <��  �
�   @  w �mD  !E  !E  =    E   j�  E  ) @E  J @�E  � "�    � '
$B  �� *	�   
 -�E  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 4E   H	F  � K�    C� N	�   "8 QR   t TR    . V�E  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   4E  sF  ! 	R hF  F  �F  ! 	� F  
K   r9I  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m H #	�I  �  '
�I   �^   (1    .�   )	�   (o�   -1   0i�   .	�   8��   /
�I  < �   �I  =    �   �I  =    �   09I  	p�  !Ls.  	t�  !M�I  	K�  !N�I  	x�  !O�I  	��  !P�I  	��  !Q�I  	r�  !R�I  �I  !J  =    	�  !SJ  	�u  !T�I  		�  !U�I  	h�  !V�I  �   aJ  =   	 	~ "8QJ  	 #V�   "  	��  $My  	(h  $N�   	l�  $N�   	�  %.y  	�  %/y  	�  %0y  	�  %2y  	w�  %8�  	�  %9�  	�  %:m  	�_  %;�   	��  %>y  	�  %Jy  	"�  %R�  	t�  %S�   	�w  %T�   	؜  %Y�   	q�  %[y  	Ƚ  %^�  	�  %_�   	�y  %`�   	b�  %c�   	+�  %fy  	��  %iy  	֘ %l�   	�J  %x�   	��  %y�   	ks  %�   	�  %��   	J�  %��   	�i  %��   	��  %�y  	��  %�y  	��  %�y  	<� %�y  	��  %�y  	��  %�y  	5�  %�y  	<m  %��   	 K  %��   	�R  %��   	op  %��   	�m  %��   	D  %��   	X�  %��   	If  %��   	� %��   	��  %�y  	�U  %�y  	`  %�y  	J�  %�y  	��  %�y  	� %��  �7  M  =    	�  %��L  y  'M  =    	� %�M    CM  =   	 	,�  %�3M  	R�  %�[M      qM  =    	�u  %�aM  	��  %�9  	�e  %��   �   �M  =   � 	(�  %��M  	�  %�y   ��  %�   �v  %�    n�  %�    4�  %�    *b %�    ��  %yJ  *�s -�   	Wf     +�?  6	 Yf     +�?  7	 Wf     +�?  8	 ^f     +	@  9	 Wf      �n P�  ,�t ��)A           �P  -m�  �~0  9� 3� -*� ��'  �� �� .th �~0  �� �� .an ��  ,� &� .x ��  x� v� .y ��  �� �� .z ��  �� �� /�  ��  � � 0�)A     �]  _O  1U| 1Tv 1Q@F$ 0*A     �]  �O  1U| 1Ts 1Q@F$ 0%*A     �]  �O  1U| 1Ts 1Q@F$ 0W*A     pW  �O  1R~  0p*A     ^  �O  1Uv  2�*A     ^  2�*A     ^  0�*A     ^  P  1T}  3�*A     �Q   4�j �~0  �(A           �LQ  -m�  �~0  �� �� -`5 �~0   � �� -*� ��'  R� L� .th �~0  �� �� .an ��  �� �� /S� �
�   /� '� 0�(A     pW  �P  1R�Q 0�(A     ^  �P  1Us  2)A     ^  2&)A     '^  2.)A     '^  2Z)A     ^  2t)A     ^  2�)A     3^  5�)A     �Q  1Us   4�e �	~0  �(A     -       ��Q  -y �!~0  �� �� 6�(A     $       7�s �f.  	 �e       ,�s �4(A     [       �R  8th �#~0  �� �� 2=(A     '^  0�(A     ?^  R  1Us  9�(A     �[  1U�U  ,cq n�'A     �       ��R  8x o�  �� }� 8y p�  �� �� 8z q�  � � -\q r�   �� y� .th t~0  � � 2�'A     '^  2�'A     '^  0�'A     pW  �R  1U�\�1Tw �1R& 2�'A     '^  3+(A     \   ,�e S'A     �       ��S  8x T�  �� �� 8y U�  �� �� 8z V�  	� � .th X~0  w� o� 2)'A     '^  20'A     '^  0J'A     pW  �S  1U�\�1T�X�1R% 2Y'A     '^  9�'A     \  1T_  ,�s �7%A     �      ��T  -cp �#[M  �� �� .i ��   m� g� .bit ��   �� �� /y �~0  �� �� .x ��  0� .� .y ��  U� S� .z ��  z� x� :�%A     �T  �T  1U�U 0&A     K^  �T  1U	h�B      2�&A     pW  2�&A     '^   , ��#A     L      ��U  -cp �![M  �� �� .p ��:  � � .x ��  -� )� .y ��  s� o� .z ��  �� �� /y �~0  �� �� .i ��   $� � 0/$A     W^  �U  1Us  0I$A     pW  �U  1Q@K$1R0 0�$A     c^  �U  1U|  2(%A     o^  31%A     {^   ,�s \�"A     2      ��V  .x ^�  �� �� .y _�  �� �� .z `�  �� �� .ss bI:  � � .mo c~0  F� @� /cp d[M  �� �� .i f�   �� �� 0##A     �^  �V  1Uv 1T|  07#A     pW  �V  1Uv 1T| 1R( 0D#A     ^  �V  1TZ 5�#A     pW  1Uv 1T|   ,11 <�A     �       �pW  -y <~0  B� :� 0=A     �^  BW  1Us  0EA     �^  ZW  1Us  9NA     �^  1U�U  4�( �~0  �A     +      �kX  8x ��  �� �� 8y ��  �� �� 8z ��  K� E� -*� ��'  �� �� /y  ~0  �� �� ;st �,  <y� z,  0�A     �^  1X  1U�1T51Q0 2A     '^  0kA     �^  VX  1Us  5�A     �^  1Us   ,ut �"A     �       �Y  -y �~0  J� 8� 0'"A     P[  �X  1Us  0N"A     �Z  �X  1Us  :t"A     \  �X  1U�U 2�"A     '^  9�"A     Y  1U�U  ,Rt � A           ��Z  -y ~0  � � .x ��  �� �� .y ��  �� �� .z ��  � � .ss �I:  =� ;� .mo �~0  h� `� /cp �[M  �� �� 0!A     �^  �Y  1Us 1Tv 1Q|  08!A     pW  �Y  1R' 0E!A     ^  	Z  1T# 0O!A     �^  'Z  1Uv 1T|  0c!A     pW  KZ  1Uv 1T| 1R' 0p!A     ^  cZ  1T# 0�!A     pW  �Z  1Uv 1T|  9�!A     �V  1U�U  =t �5A     �      �P[  >mo �~0  +� � ?S� ��  �� �� ?� ��  �� �� @p  B[  /�s 1�   �� �� 0"A     ^  ,[  1Us 1T" 9ZA     �[  1U�U  2�A     3^   A4t l�[  Bmo l~0  C�s n�  C�t o�  C�R  p�:  C�p q�  C	q r�   =�s T�A     m       �\  >mo T ~0  �� �� 0�A     \  �[  1Us  2�A     '^  93A     ^  1U�U  D�e 0y  NA     z       ��\  Ey 1~0  �� �� E�� 2�#  �� �� Fst 4�,  @� <� 0kA     �V  �\  1Us  G�A     1Us   HP[  �A     5      ��]  I][  �� x� Jh[  Jt[  J�[  J�[  J�[  KP[  �  �]  I][  Z� N� L�  Mh[  �� �� Mt[   � � M�[  Z� V� M�[  �� �� M�[  +� � 0�A     ?^  P]  1Us  0�A     �^  h]  1Us  :�A     �V  �]  1U�U 0�A     �[  �]  1Us  0� A     \  �]  1T� 0� A     ^  �]  1T
 � 5� A     ^  1T
 �   9�A     \  1U�U  Ncg cg �N� � #6Nd  d  "	NEf Ef xN� � &!N�h �h �	N\i \i �	N��  ��  '7N�- �- %Net et NNt t !1N�4 �4 "/N3, 3, �Ni i �N(t (t #9Nc c HN� � 6N�d �d �N3b 3b GN�" �" �	N�q �q � �P   �z  S#  �t �*  �*A     �      	� r�  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �   	"  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�  4  
K   "z  ��  WH  �~  �O  �m  ��   �  ��  ��  	 
K   	�  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  	(z  
K   	/�  ��   [r  �4 #�  �   �X  	5�  
K   	:m  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  	K
  
�   	P�  =_  ��   R�  N�  ��  ��   �p  	Wy  
K   
3�  ��   ({  ��  ğ   F]  
8�  
K   
Y$  ��   �c  |  ��  l  ��  �   
K   
ku  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  
{$  
K   
��  &�   �  º  GY  �f  ��   v�  
��  
K   
��  GQ   ϼ  �  �_  X  &�  �b   t�   �   �      =   �' 
  	��  1  	]  48      O  =   � >  	Zy  8O  �  v  =   =   � `  	��  ;v  Ʃ  QK   �  �  �  =     �  	�  W�  �p  #�  �  �   S�  $�  �  �  R    T}  %�      R   R    '	@  acv )�  ��  *�  ��  +�   �y -  �Y  6@  ��  :�  s�  <�   �H  =�  xz  >L   X  x @X  B  �  =    4  �  =    
�	  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x ��  
K   c
  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �  
K   ��#  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  uo
  (x	p$  �u zc
   � {	�   s |	�   � ~@  N�  �#  ��  �	�   ��  �	�     J]  �$  p$  �$  =   �  �^  �}$  �   �$  !  �  ��$  "K   ��'  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �$  \	Y)  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /(  Y)  v)  =   �  ��  1f)  �]  ��Y+  `e ��   x ��  y ��  z ��   ��  �Y+  (cN  �Y+  0Mp ��  8�u �c
  <� ��   @�H  �Y+  Hr�  �Y+  P��  ��+  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� ��'  �y� ��+  �s ��   ��� ��+  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  Y+  ���  �   ���  	�   ��R  �-  �f�  �   �I}    ���  Y+  � �)  Gx  ��+  >} ��0   �}  �B  �|  �B  
 _+  Y)  p$  #d  HN�-  mo P�/   ��  Q�6  cmd R"  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g�6  8�W  h�6  P��  iy  h�� l�/  l�N  mu  |E�  pu  ��W  r�6  �~�  s�/  �*� t�/  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��/  �$�R  ��    $��  ��   $�  ��   $h  ��6  $I�  �y  @ �+  �z �)  �  	��  ��   	�\  �y  	�  ��-  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  ��-  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	t.  x E�   y F�   �{ HT.  (T	�.  `e V�   x W�  y X�  z Y�    	�  [�.  �a	�/  = c�   F�  d�  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  o�/  ��  r
�/   iK  u�.  0��  x
�   XS�  {�/  `��  ~R   h��  ��   pu| �t0  x �-  �   �/  =    �}  X�t0  v1 �)1   v2 �)1  dx ��  dy ��  �  �B  �k �B  tag �B  �W  ��  �o �/1  $��  �1  4SX  ��0  8d�  ��0  @��  �
�   H��  �R   P z0  �/  �z ��.  �	�0  2�  ��   ]  ��  �h  �B  �N  �B  
�K  �B  >} ��0   �0  �}  ��0  
K   �1  ��   �  o�  ��   ��  ��0  t.  �  ?1  =    �u  ��/  �z �_+  8�	�1  v1 �)1   v2 �)1  82  ��  Mp ��  [�  ��1   �  ��1   SX  ��0  (d�  ��0  0 �0  ?1  A{ �W1  4	82  %x �   %y 	�  %dx 
�  %dy �  �o 82  )�  �  0 �  N2  =   =    (} �1  �  *�  &v  @23  @�  43   %x1 5�   %x2 6�   .]  8�  5]  9�  �� :�  ��  =�   �  @�   ��  C�  $�n  G#3  (9x  H#3  0�^  I#3  8 �1  B  >�  Kh2  &�h  PR4  s�  U4   �H  V4  %x1 X�   %x2 Y�   %gx \�  %gy ]�  %gz `�   %gzt a�  $�x  d�  (� f�  ,~�  i�  0t  k�  4.� l�   8�  p4  @	�  r�   H 63  [2  �h  t63  �	`4  �c  �y   �O  �`4  �x  �
p4   B  p4  =    �  �4  =    I�  �+4  �	�4  �  ��    �  ��4   �4  �  ��4  '��	q5    ��   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  %top �	q5  (��  �	�  U(��  �	�  V(� �	q5  W(�  �	�  � �  �5  =   ? ��  ��4  	�5  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�5  �5  6  =    	S�  '�5  
K   706  {�   U�  ~�   >	l6  �� @�+   s A
�   sx B�  sy C�   Nz E06  
K   1�6  ��   ��  ��   �y  9x6  �   �6  =    y  �6  =    y  �6  =    l6  �6  =    hy ��+  (�	U7  in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�/  �a  �
�   $ ��  ��6  ��	�7  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��7  ( U7  
8  =    ޴  �a7  	.L  &"8  �  	׮  )"8  	�  +"8  	�  ,"8  	�Q  .4  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�8  �   	��  8�8  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�8  �4  	��  H�   	��  I)1  	��  K�   	a� L3  	w�  N�   	P{ O�0  	��  Q�   	��  RH9  K1  	��  T�   	�� Uf9  N2  	�}  W�   	u| X�1  	M�  Z�   	P�  [�1  	��  a�  	��  b�  	�  c�  	�p  e�  	�T  f�9  �6  	�a  j�  �   �9  =   � 	ը  l�9  �  :  =   @ 	�p  m:  	 �  p�  	p|  q�  	$Y  v�   	�K  y�   	g  {`:  �5  	d�  |`:  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   4  ;  =   =   / 	��  E;  4  4;  =   / 	Ԁ  F$;  4  V;  =   =    	7� G@;  	�R  I�   	��  J4  	��  U�   	P�  \.  	��  ].  	L�  ^.  	ߵ  _.  	�  a.  	@�  3  	[�  �1  	 �  �1  	SX  �0  	d�  �0  	��  �   	_�   �   	��  "y  	��  %y  	'�  &y  	�]  (y  )3  V<  =   � 	�P  *F<  	ӯ  +n<  )3  	|  -�<  4  	��  .�<  	��  /�<  �<  �<  �   �    	��  #3  �   �<  	qY  "�<  	�  #�<  B  �<  =   ? 	��  %�<  	��  &�<  �  =  =   � 	@Y  (=  �  :=  =   ? 	V�  ))=  4  V=  =    	�h  F=  	�  n=  4  	�  4  	�f  !�<  	r�  "�<  	��  %#3  	��  &#3  	׆  '�  	��  (�  	�  *�  	��  +�  	�  4  	��  �   	�_  �   	�_  �   	b  �  	t  �  	j�  "�-  	�  :�   	��  ;�   	��  <�   	�W  >4  	hn  @�  	U~  A�  	�  B�  	 �  C�  	%�  F�-  	�u  H�-  	z  I�-  	ʓ  C�    �>  =    	��  b�>  �   �>  =    	��  c�>  	0K  d�   	?�  e�   �	L?  x ��   y ��  dx ��  dy ��   ��  �?  �z?  �p �
�/  ��  �
�1   �	�?  {q ��   ��  �y  d �	X?   t�  �z?  �?  �?  =   � 	r ��?  	�T  ��?  �?  	l�  ��  	�  ��  	?k  ��  	�d  ��  	2~ �L?  	��  �y  	��  ��  	k�  ��  	Z�  ��1  �1  _@  =    	�v  �O@  	�v  ��   	"�  ��/   �  �-   �U  #3   ��  #3   t�  �    �  	�    .Y  
�   7Y  �   �h  �@  �/   *� �/   <i  �/  	G  y  	��  �   �   3A  =    
K   �TA  )top  �G  �  �]  �3A   �	�A  ��  ��1   ��  �TA  O{  �
�   ��  �
�   iK  ��A   �.  ��  �`A  �A  �A  =    	��  ��A  "K    B  )up  �  �F  �S   FT  
�A  "K   ;B  ��   �x  H�  ��  �H   ��  B  H	�B  `e �   >} �0  L� �   %low �  $+�  �  (�Z !
�   ,r� "
�   0�f  # B  4�f  $ B  8��  %y  <%tag &
�   @*� ';B  D �w )HB  C  C  =    �B   �  2C  "K   �_C  ��   �s  z�  ��  �T  ܭ   gY  �+C  H�	D  `e ��   *� �_C  >} ��0   �W  ��  (�}  ��  ,L� ��  0��  �y  4��  �
�   8%tag �
�   <��  �
�   @  w �lC   D   D  =    D   j�  D  "K   XTD  )ok  �b �b  Mb ]3D  ) mD  J @�D  � "�    � '
#A  �� *	�   
 -�D  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 aD   H	AE  � K�    C� N	�   "8 QR   t TR    . VE  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   aD  �E  ! 	R �E  AE  �E  ! 	� �E  
K   rfH  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	  V�   "  	��  !My  	(h  !N�   	l�  !N�   	�  ".y  	�  "/y  	�  "0y  	�  "2y  	w�  "8�  	�  "9�  	�  ":m  	�_  ";�   	��  ">y  	�  "Jy  	"�  "R�  	t�  "S�   	�w  "T�   	؜  "Y�   	q�  "[y  	Ƚ  "^�  	�  "_�   	�y  "`�   	b�  "c�   	+�  "fy  	��  "iy  	֘ "l�   	�J  "x�   	��  "y�   	ks  "�   	�  "��   	J�  "��   	�i  "��   	��  "�y  	��  "�y  	��  "�y  	<� "�y  	��  "�y  	��  "�y  	5�  "�y  	<m  "��   	 K  "��   	�R  "��   	op  "��   	�m  "��   	D  "��   	X�  "��   	If  "��   	� "��   	��  "�y  	�U  "�y  	`  "�y  	J�  "�y  	��  "�y  	� "��  �6  K  =    	�  "��J  y   K  =    	� "�K    <K  =   	 	,�  "�,K  	R�  "�TK      jK  =    	�u  "�ZK  	��  "�
8  	�e  "��   �   �K  =   � 	(�  "��K  	�  "�y   ��  "�   �v  "�    n�  "�    4�  "�    *b "�    ��  "rH  *C  &
	@^f     +�t #X-A     E       ��L  ,+w #!C  �� �� -i %
�   "� � .y-A     P  wL  /U�U 0�-A     P  /U	��B       +�t E+A     -       ��L  ,+w C  �� �� -i 
�   �� �� 0r+A     P  /U	��B       +�t 	+A     <       �8M  1��  �1  U-j 	
�   +� %�  2�t ��*A     2       �wM  3tag ��   U4i �
�   }� w�  5�t ��   r+A     �      �(O  6��  ��1  �� �� 6*� �;B  !� � 6�m ��   s� m� 7+w �C  �� �� 7�k �
�   � � 4rtn �
�   �� �� 4sec ��0  � � .�+A     8M  =N  /Uu  .�+A     P  [N  /Uv /T}  .�+A     %P  }N  /UH/T6/Q0 .�+A     1P  �N  /Us  .W,A     =P  �N  /U  .�,A     IP  �N  /U  .�,A     IP  �N  /U  .-A     UP  �N  /U  8"-A     aP  .5-A     mP  O  /U|  8B-A     �L   2�t -�-A     .      �P  6+w -C  c� S� 4res /TD      .�-A     yP  �O  /X0/Y1 ..A     mP  �O  /TF .Q.A     mP  �O  /TC 9f.A     L  �O  /U�U .~.A     yP  �O  /R0/X0/Y	� :�.A     mP   ;c c H;��  ��  #7;Vb Vb `;� � 6;3b 3b G;�k �k X;l l T	;Nk Nk U	;� � $!;� �  6<c c ` e`    ~  S#  �u �*  �.A     �      ?� #�  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �  
K   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
K   /  ��   [r  �4 #�  �   �X  5�  
K   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K&  
�   P�  =_  ��   R�  N�  ��  ��   �p  W�  
K   3�  ��   ({  ��  ğ   F]  8�  
K   Y@  ��   �c  |  ��  l  ��  �   
K   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {@  
K   ��  &�   �  º  GY  �f  ��   v�  ��  
K   �  GQ   ϼ  �  �_  X  &�  �b   
K   	Kf  � � ^�  �� e  2 8� ��  �  _�  �   t�  
 �   f  r  �  =   �' w  	��  1�  	]  4�  r  r  �  =   � �  	Zy  8�  �  �  =   =   � �  	��  ;�  Ʃ  QK   �       =       	�  W  �p  #3  9  @   S�  $L  R  ]  R    T}  %i  o    R   R    '	�  acv )'  ��  *@  ��  +]   �y -  �Y  6�  ��  :�  s�  <�   �H  =�  xz  >�   �  x @�  B    =    4  ,  =    
�	s  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x �,  
K   �	  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �  
K   �c#  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�	  (x	�#  �u z�	   � {	�   s |	�   � ~�  N�  c#  ��  �	�   ��  �	�     J]  �p#  �#  �#  =   � �^  ��#  �   $    �  �$  !K   �l'  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o   $  \	�(  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /y'  �(  �(  =   � ��  1�(  
K   p�)  �! 9& +! v( %# 0  B& @�! ��"  w#  	$  �-  S%  �)   0  @&  ��"    !0    m0    b-    �.    �$     /   @ %   � <"    U-    5'    	!  �]  ���+  `e �    x �f  y �f  z �f   ��  ��+  (cN  ��+  0Mp ��  8�u ��	  <� ��   @�H  ��+  Hr�  ��+  P��  ��+  X��  �f  `m�  �f  d��  �f  h  �f  l3F  �f  p8F  �f  t=F  �f  x��  ��   |*� �l'  �y� ��+  �s ��   ��� ��+  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  �+  ���  �   ���  	�   ��R  �-  �f�  �   �I}  s  ���  �+  � �)  Gx  ��+  >} �11   �}  �B  �|  �B  
 �+  �(  �#  "d  HN�-  mo P�/   ��  Q~7  cmd RQ7  �  Wf  (_  Yf   #_  [f  $bob ]f  (�  a�   ,�[  b�   0sb  d�   4d]  g�7  8�W  h�7  P��  iy  h�� l�/  l�N  m�  |E�  p�  ��W  r�7  �~�  s�/  �*� t�/  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��/  �#�R  ��    #��  ��   #�  ��   #h  ��7  #I�  �y  @ �+  �z �)  �  	��  ��   	�\  �y  	�  �
.  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  ��-  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	�.  x Ef   y Ff   �{ H�.  (T	/  `e V    x Wf  y Xf  z Yf    	�  [�.  �a	�/  = cf   F�  df  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  o�/  ��  r
�/   iK  u/  0��  x
�   XS�  {�/  `��  ~R   h��  ��   pu| ��0  x �-  �   0  =    �}  X��0  v1 �v1   v2 �v1  dx �f  dy �f  �  �B  �k �B  tag �B  �W  �  �o �|1  $��  �j1  4SX  �11  8d�  �11  @��  �
�   H��  �R   P �0  0  �z �/  �	11  2�  �f   ]  �f  �h  �B  �N  �B  
�K  �B  >} �11   �0  �}  ��0  
K   �j1  ��   �  o�  ��   ��  �C1  �.  f  �1  =    �u  �0  �z ��+  8�	2  v1 �v1   v2 �v1  82  �f  Mp ��  [�  �2   �  �2   SX  �11  (d�  �11  0 71  �1  A{ ��1  4	�2  $x f   $y 	f  $dx 
f  $dy f  �o �2  )�    0 f  �2  =   =    (} ,2  �  *�  %v  @2j3  @�  4j3   $x1 5�   $x2 6�   .]  8f  5]  9f  �� :f  ��  =�   �  @f   ��  Cf  $�n  Gp3  (9x  Hp3  0�^  Ip3  8  2  B  >�  K�2  %�h  PR_4  s�  U_4   �H  V_4  $x1 X�   $x2 Y�   $gx \f  $gy ]f  $gz `f   $gzt af  $�x  df  (� ff  ,~�  if  0t  kf  4.� l�   8�  pe4  @	�  r�   H �3  �2  �h  t�3  �	�4  �c  �y   �O  ��4  �x  �
�4   B  �4  =    �  �4  =    I�  �x4  �	5  �  ��    �  �5   �4  �  ��4  &��	�5    �f   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  $top �	�5  '��  �	�  U'��  �	�  V'� �	�5  W'�  �	�  � �  �5  =   ? ��  �5  	46  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�5  46  P6  =    	S�  '@6  
K   7}6  {�   U�  ~�   >	�6  �� @�+   s A
�   sx Bf  sy Cf   Nz E}6   	Q7  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�6  
K   1~7  ��   ��  ��   �y  9]7  �   �7  =    y  �7  =    y  �7  =    �6  �7  =    hy ��+  (�	:8  in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�/  �a  �
�   $ ��  ��7  ��	�8  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��8  ( :8  �8  =    ޴  �F8  	.L  &9  f  	׮  )9  	�  +9  	�  ,9  	�Q  .e4  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7y9  �   	��  8y9  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�9  5  	��  H�   	��  Iv1  	��  K�   	a� Lj3  	w�  N�   	P{ O11  	��  Q�   	��  R-:  �1  	��  T�   	�� UK:  �2  	�}  W�   	u| X2  	M�  Z�   	P�  [2  	��  af  	��  bf  	�  cf  	�p  e�  	�T  f�:  �7  	�a  j�  �   �:  =   � 	ը  l�:  �  �:  =   @ 	�p  m�:  	 �  pf  	p|  q�  	$Y  v�   	�K  y�   	g  {E;  �5  	d�  |E;  	��   f  		�  !f  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +f  	`�  ,f  	A�  -f  	��  /�   	��  1�   	P�  2�   e4  �;  =   =   / 	��  E�;  e4  <  =   / 	Ԁ  F	<  e4  ;<  =   =    	7� G%<  	�R  I�   	��  Je4  	��  U�   (	P�  \x<  k<  	��  ]x<  	L�  ^x<  	ߵ  _x<  	�  ax<  	@�  j3  	[�  2  	 �  2  	SX  11  	d�  11  	��  �   	_�   �   	��  "y  	��  %y  	'�  &y  	�]  (y  v3  B=  =   � 	�P  *2=  	ӯ  +Z=  v3  	|  -l=  e4  	��  .l=  	��  /l=  �=  �=  �   �    	��  p3  �   �=  	qY  "�=  	�  #�=  B  �=  =   ? 	��  %�=  	��  &�=  f  	>  =   � 	@Y  (�=  f  &>  =   ? 	V�  )>  k4  B>  =    	�h  2>  	�  Z>  k4  	�  k4  	�f  !�=  	r�  "�=  	��  %p3  	��  &p3  	׆  'f  	��  (f  	�  *f  	��  +f  	�  e4  	��  �   	�_  �   	�_  �   	b  f  	t  f  	j�  "�-  	�  :�   	��  ;�   	��  <�   	�W  >e4  	hn  @f  	U~  Af  	�  Bf  	 �  Cf  	%�  F�-  	�u  H�-  	z  I�-  	ʓ  C   s  �?  =    	��  b�?  �   �?  =    	��  c�?  	0K  d�   	?�  e�   �	8@  x �f   y �f  dx �f  dy �f   ��  � @  �f@  �p �
�/  ��  �
2   �	�@  {q �f   ��  �y  d �	D@   t�  �f@  �@  �@  =   � 	r ��@  	�T  ��@  �@  	l�  �f  	�  �f  	?k  �f  	�d  �f  	2~ �8@  	��  �y  	��  �f  	k�  �f  	Z�  �2  2  KA  =    	�v  �;A  	�v  ��   	"�  ��/  �  �-  �U  p3  ��  p3  t�  �   �  	�   .Y  
f  7Y  f  �h  �A  �/  *� �/  <i  �/  	G  y  	��  �   �   B  =    
K   �@B  )top  �G  �  �]  �B   �	�B  ��  �2   ��  �@B  O{  �
�   ��  �
�   iK  ��B   /  ��  �LB  �B  �B  =    	��  ��B  !K   �B  )up  �  �F  �S   FT  
�B  !K   'C  ��   �x  H�  ��  �H   ��  �B  H	�C  `e     >} 11  L� f   $low f  $+�  f  (�Z !
�   ,r� "
�   0�f  #�B  4�f  $�B  8��  %y  <$tag &
�   @*� ''C  D �w )4C  D  D  =    �C  �  2�C  !K   �KD  ��   �s  z�  ��  �T  ܭ   gY  �D  H�	�D  `e �    *� �KD  >} �11   �W  �f  (�}  �f  ,L� �f  0��  �y  4��  �
�   8$tag �
�   <��  �
�   @  w �XD  E  E  =    �D  j�  �D  ) +E  J @�E  � "�    � '
B  �� *	�   
 -�E  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 E   H	�E  � K�    C� N	�   "8 QR   t TR    . V�E  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   E  ^F    	R SF  �E  uF    	� jF  
K   r$I  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	  V�   Q7  	��  !My  	(h  !N�   	l�  !N�   	�  ".y  	�  "/y  	�  "0y  	�  "2y  	w�  "8  	�  "9�  	�  ":�  	�_  ";�   	��  ">y  	�  "Jy  	"�  "R�  	t�  "S�   	�w  "T�   	؜  "Y�   	q�  "[y  	Ƚ  "^�  	�  "_�   	�y  "`�   	b�  "c�   	+�  "fy  	��  "iy  	֘ "l�   	�J  "x�   	��  "y�   	ks  "�   	�  "��   	J�  "��   	�i  "��   	��  "�y  	��  "�y  	��  "�y  	<� "�y  	��  "�y  	��  "�y  	5�  "�y  	<m  "��   	 K  "��   	�R  "��   	op  "��   	�m  "��   	D  "��   	X�  "��   	If  "��   	� "��   	��  "�y  	�U  "�y  	`  "�y  	J�  "�y  	��  "�y  	� "��  �7  �K  =    	�  "��K  y  �K  =    	� "��K  s  �K  =   	 	,�  "��K  	R�  "�L  s  s  (L  =    	�u  "�L  	��  "��8  	�e  "��   �   ]L  =   � 	(�  "�LL  	�  "�y  ��  "�  �v  "�   n�  "�   4�  "�   *b "�   ��  "0I  *v d
f  	4_f     *�u e
f  	8_f     + s _
f  	0_f     ,�u \:A     [       ��M  -�R  \ �:  i  c  .i ^
�   �  �  .psp _�M    /�� `�+  o m 0V:A     +^  1Us 1Tv   �6  ,et H�9A     $       ��M  -�R  H!�:  � � .i J	�   � � 2:A     F]  1U�U  ,%u ;�9A            �RN  -�R  <�:  % ! 3psp =�M  b ^ 2�9A     �_  1T9  ,�v N9A     �       �'O  3mo �/  � � .i �   � � .j �     /\q �   r n .an �  � � 4u9A     �_  �N  1Q@F$ 4�9A     �_  O  1R* 5�9A     `  0�9A     `  1R|   ,Fu C9A            �eO  6�R  �:  U7psp ,�M  T ,=u 89A            ��O  6�R  �:  U7psp ,�M  T ,�v -9A            ��O  6�R  �:  U7psp ,�M  T ,(v �x8A     �       ��P  -�R  ��:  � � 3psp ��M  w m 4�8A     �_  AP  1T1 4�8A      `  YP  1T� 4�8A     �V  wP  1Us 1Qq  4	9A     +^  �P  1T1 59A     mT  8)9A     �S   ,Qv ��7A     �       �R  -�R  ��:  � � 3psp ��M  B > .i �
�   � { /Mp ��  � � /\q �
�     4�7A     �_  FQ  1T4 4�7A      `  ^Q  1T� 4�7A     �V  |Q  1Us 1Qq  48A     +^  �Q  1T1 5	8A     mT  58A     `  58A     `  5$8A     `  5+8A     `  598A     `  0g8A     ,`  1Tv 1Q@G$1X } #5  ,Cv �,7A     p       ��R  -�R  ��:  h b 3psp ��M  � � .i �
�   � � 4D7A     �_  �R  1T2 4Q7A      `  �R  1T� 4k7A     �V  �R  1Us 1Qq  4�7A     +^  �R  1T1 5�7A     mT  0�7A     �S  1T0  ,u ��6A     m       ��S  -�R  ��:  R L 3psp ��M  � � 4�6A     �_  OS  1T1 4�6A      `  gS  1T� 4�6A     �V  �S  1Us 1Qq  47A     +^  �S  1T1 57A     mT  8,7A     �S   ,u {Z6A     e       �mT  3mo |�/  � � -v }y  H B /Mp �  � � /\q �
�   � � 5l6A     `  5�6A     `  5�6A     `  2�6A     ,`  1U�U1Q@G$  , u b�5A     e       �&U  3mo b�/  	 		 .an d�  i	 [	 4
6A     �_  �T  1Uv 1Ts 1Q@F$ 4-6A     �_  U  1Uv 1Ts��� 1Q@F$ 0P6A     �_  1Uv 1Ts���`1Q@F$  ,0u K�5A     R       ��U  -�R  L�:  
 
 3psp M�M  h
 d
 4�5A     �V  �U  1Uu 1Qq  5�5A     `  4�5A     +^  �U  1Us 1T1 2�5A     8`  1T"  ,Wu <}5A     &       �HV  -�R  =�:  �
 �
 3psp >�M  �
 �
 4�5A     �V  3V  1Uu 1Qq  2�5A     8`  1T#  ,�u /W5A     &       ��V  -�R  0�:    3psp 1�M  \ X 4o5A     �V  �V  1Uu 1Qq  2}5A     8`  1T!  9�u �.A            �W  6�R  $�:  U6iv 0�   T6�m =�   Q ,v �\4A     �       �NX  -�R  ��:  � � 3psp ��M    /Mp ��  _ Q /\q �
�    � /�  �
�   u q 5k4A     `  5{4A     `  5�4A     `  4�4A     �_  �W  1Ts 1Q @  4�4A     ,`  X  1Ts 1Q @ 1X| :1$# :�4A     �_  )X  1T< 4�4A     �_  @X  1T= 55A     D`   ,Ou ��3A     �       �iY  -�R  ��:  � � 3psp ��M   � /Mp ��  > : /\q �
�   x t /�  �
�   � � 5�3A     `  5�3A     `  5�3A     `  44A     �_  Y  1Ts 1Q@B$ 44A     ,`  CY  1Ts 1Q@B$1X�\� 444A     �_  [Y  1TS 5P4A     D`   ,�v ��3A     ,       ��Y  -�R  ��:  � � 3psp ��M  ? ; 4�3A      `  �Y  1T� 2�3A     +^  1U�U1T1  ,�v �S3A     .       �VZ  -�R  ��:  | x 3psp ��M  � � ;`v �c#  2�3A     +^  1U�U1T0  ,�v x3A     >       ��Z  -�R  y�:  � � 3psp z�M  { q :D3A     +^  �Z  1U�U1T01Q0 2R3A     F]  1U�U  ,�u e3A            �7[  -�R  f�:  � � 3psp g�M  1 - 23A     ]  1U�U  ,�h N�2A     /       ��[  -�R  O�:  r j 3psp P�M  � � :3A     �\  �[  1U�U 23A     ]  1U�U  ,au �1A            ��\  -�R  �:  P > 3psp �M  "  ;`v c#  /Mp 
�   � � 42A      `  2\  1T� 4,2A     �_  I\  1T; :V2A     +^  g\  1U�U1T0 :�2A     �\  �\  1U�U 5�2A     P`  5�2A     P`   ,Nl  �1A            ��\  -�R   �:  
  2�1A     +^  1U�U1T0  <�v �]  =�R  ��:  >`v �c#   ?�u �	y  F]  =�R  � �:  >~�  ��  >r� ��    @3v ��/A     [       ��]  A�R  �!�:  K C B`v �c#  � � 4 0A     �_  �]  1T: 2/0A     +^  1U�U1T0  @ v g�/A     M       �+^  A�R  g�:  � � B"v if    >Mp j
�   5�/A     P`  5�/A     P`   @�u 2�.A     �       ��^  A�R  3�:  8 2 A@�  4�   � � A 5c#  � � Cpsp 7�M    B�� 8�+  b \ Dt/A     1Uv 1T|   E]  /0A     _      �9_  F!]  � � G-]    G9]  ? ; H]  �  I!]  J�  K-]  K9]  0�1A     +^  1T0    E�\  �1A     ?       ��_  F�\   u K]  L�\     �_  F�\  � � J   K]  4�1A      `  �_  1T� 4�1A     +^  �_  1Us 1T0 8�1A     \`    0�1A     ]  1Us   M� �  6Mcg cg �M�( �( kM� � #!Ndj dj M�e �e s	Mf f �M�t �t yMEf Ef xMd  d  
"	MWj Wj  �y   m�  S#  zw �*  t:A     �      ռ �  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  9�  
�   3   	Y�  %(  	��  &(  0t  W  e2    �0  }  �x �D   ��  K  �� 0s  K   J�  D   �C  
D  ���� �C  N�  ڵ  R  �  	"|  *�  	��  +�  	I�  ,�  	�a  -�  	 	�  ��  	"e   E�  	#e  e% 	$l  u  	%
�  �8 	&
�  ��  	)
�  /b  	-
�  ��  	.	�   a  	2
�  �T  	3
�   Mx 	4  �  K   
"�  ��  WH  �~  �O  �m  ��   �  ��  ��  	 t�   �   �  
�    =   �' �  	��  1  	]  4+  �  
�  B  =   � 1  	Zy  8B  
�  i  =   =   � S  	��  ;i  Ʃ  QK   z  
�  �  =     �  	�  W�  K   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  K   /1  ��   [r  �4 #�  �   �X  5  K   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K=  �   P�  =_  ��   R�  N�  ��  ��   �p  W�  K   3  ��   ({  ��  ğ   F]  8�  K   YW  ��   �c  |  ��  l  ��  �   K   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {W  K   ��  &�   �  º  GY  �f  ��   v�  ��  K   �,  GQ   ϼ  �  �_  X  &�  �b   �p  #8  >  E   S�  $Q  W  b  R    T}  %n  t  �  R   R    '	�  acv ),  ��  *E  ��  +b   �y -�  �Y  6�  ��  :�  s�  <�   �H  =�  xz  >�   �  x @�  
l  !  =    
^  1  =    
�	x  x �l   y �l  Mp �l  *� �l  ޽  �l   ~x �1  K   �
  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  K   �h$  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�
  (x	�$   �u z�
    � {	�    s |	�    � ~�   N�  h$   ��  �	�    ��  �	�     J]  �u$  
�$   %  =   � !�^  ��$  !�  �(  "K   �f(  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  %  \	�)   �Y  	�     *O  	�    ��  	�    �  	�    b�  	�    ��  	�    �  	�    +�  	�    Zp  	�     o�   	�   $ m�  !	�   ( 4�  "	�   , �  #	�   0 �  $	�   4 ��  %	�   8 L� &	�   < ��  '	�   @   (	�   D ��  )	�   H \q *	�   L z�  +	�   P �  ,	�   T /�  -	�   X ʤ  /s(  
�)  �)  =   � !��  1�)  �]  ���+  `e �   x ��  y ��  z ��   ��  ��+  (cN  ��+  0Mp �z  8�u ��
  <� ��   @�H  ��+  Hr�  ��+  P��  ��+  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� �f(  �y� �,  �s ��   ��� �,  ��  ��   ��  ��   �ʺ  ��   ��l  ��   �  �  �+  � ��  �   � ��  	�   � �R  �-  � f�  �   � I}  x  � ��  �+  � �)  Gx  ��+  >} �K1   �}  �l  �|  �l  
 �+  �)  �$  #d  HN�-  mo P0   ��  Q 7  cmd R�  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g7  8�W  h7  P��  i�  h�� l0  l�N  m�  |E�  p�  ��W  r,7  �~�  s0  �*� t0  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �0  �$�R  ��    $��  ��   $�  ��   $h  �<7  $I�  ��  @ ,  �z �)  �  	��  ��   	�\  ��  	�  �$.  �  	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  ��-  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	�.  x E�   y F�   �{ H�.  (T	/  `e V   x W�  y X�  z Y�    	�  [�.  �a	0  = c�   F�  d�  �~ el  h�  fl  
t�  gl  �k hl  tag il  �N  l
�   ��  o0  ��  r
0   iK  u/  0��  x
�   XS�  {0  `��  ~R   h��  ��   pu| ��0  x �-  
�   0  =    �}  X��0  v1 ��1   v2 ��1  dx ��  dy ��  �  �l  �k �l  tag �l  �W  �  �o ��1  $��  ��1  4SX  �K1  8d�  �K1  @��  �
�   H��  �R   P �0  0  �z �+/  �	K1  2�  ��   ]  ��  �h  �l  �N  �l  
�K  �l  >} �K1   �0  �}  ��0  K   ��1  ��   �  o�  ��   ��  �]1  �.  
�  �1  =    �u  �0  �z ��+  8�	.2  v1 ��1   v2 ��1  82  ��  Mp �z  [�  �.2   �  �42   SX  �K1  (d�  �K1  0 Q1  �1  A{ ��1  4	�2  %x �   %y 	�  %dx 
�  %dy �   �o �2   )�  !  0 
�  �2  =   =    (} F2  �  *�  &v  @2�3   @�  4�3   %x1 5�   %x2 6�    .]  8�   5]  9�   �� :�   ��  =�    �  @�    ��  C�  $ �n  G�3  ( 9x  H�3  0 �^  I�3  8 :2  l  >�  K�2  &�h  PRy4   s�  Uy4    �H  Vy4  %x1 X�   %x2 Y�   %gx \�  %gy ]�  %gz `�   %gzt a�  $ �x  d�  ( � f�  , ~�  i�  0 t  k�  4 .� l�   8 �  p4  @ 	�  r�   H �3  �2  �h  t�3  �	�4   �c  ��    �O  ��4   �x  �
�4   
l  �4  =    
�  �4  =    I�  ��4  �	5   �  ��     �  �5   �4  �  ��4  '��	�5     ��    �  �	�    t�  �	�    ��  �	�    /�  �	�    �  �	�  %top �	�5  (��  �	�  U(��  �	�  V(� �	�5  W(�  �	�  � 
�  �5  =   ? ��  �.5  	N6  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�5  
N6  j6  =    	S�  'Z6  K   7�6  {�   U�  ~�   >	�6  �� @,   s A
�   sx B�  sy C�   Nz E�6  K   1 7  ��   ��  ��   �y  9�6  
�   7  =    
�  ,7  =    
�  <7  =    
�6  L7  =    hy �,  (�	�7  in ��   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
0  �a  �
�   $ ��  �X7  ��	a8  2�  �
�    I�  ��  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  �a8  ( 
�7  q8  =    ޴  ��7  	.L  &�8  �  	׮  )�8  	�  +�8  	�  ,�8  	�Q  .4  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�8  �   	��  8�8  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u FI9  !5  	��  H�   	��  I�1  	��  K�   	a� L�3  	w�  N�   	P{ OK1  	��  Q�   	��  R�9  �1  	��  T�   	�� U�9  �2  	�}  W�   	u| X42  	M�  Z�   	P�  [.2  	��  a�  	��  b�  	�  c�  	�p  ez  	�T  f?:  L7  	�a  jz  
�   b:  =   � 	ը  lQ:  
z  :  =   @ 	�p  mn:  	 �  p�  	p|  qz  	$Y  v�   	�K  y�   	g  {�:  �5  	d�  |�:  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   
4  ;  =   =   / 	��  Ei;  
4  �;  =   / 	Ԁ  F�;  
4  �;  =   =    	7� G�;  	�R  I�   	��  J4  	��  U�   	P�  \�  	��  ]�  	L�  ^�  	ߵ  _�  	�  a�  	@�  �3  	[�  .2  	 �  42  	SX  K1  	d�  K1  	��  �   	_�   �   	��  "�  	��  %�  	'�  &�  	�]  (�  
�3  �<  =   � 	�P  *�<  	ӯ  +�<  �3  	|  -�<  4  	��  .�<  	��  /�<  =  =  �   �    	��  �3  �   =  	qY  "'=  	�  #'=  
l  \=  =   ? 	��  %K=  	��  &K=  
�  �=  =   � 	@Y  (t=  
�  �=  =   ? 	V�  )�=  
�4  �=  =    	�h  �=  	�  �=  �4  	�  �4  	�f  !K=  	r�  "K=  	��  %�3  	��  &�3  	׆  '�  	��  (�  	�  *�  	��  +�  	�  4  	��  �   	�_  �   	�_  �   	b  �  	t  �  	j�  "�-  	�  :�   	��  ;�   	��  <�   	�W  >4  	hn  @�  	U~  A�  	�  B�  	 �  C�  	%�  F�-  	�u  H�-  	z  I�-  	ʓ  C  
x  ;?  =    	��  b+?  
�   W?  =    	��  cG?  	0K  d�   	?�  e�   �	�?  x ��   y ��  dx ��  dy ��   ��  �{?  ��?  �p �
0  ��  �
42   �	@  {q ��   ��  ��  d �	�?   t�  ��?  
@  ,@  =   � 	r �@  	�T  �D@  @  	l�  ��  	�  ��  	?k  ��  	�d  ��  	2~ ��?  	��  ��  	��  ��  	k�  ��  	Z�  �42  
42  �@  =    	�v  ��@  	�v  ��   	"�  �0  !�  �-  !�U  �3  !��  �3  !t�  �   !�  	�   !.Y  
�  !7Y  �  !�h  RA  0  !*� 0  !<i  0  	G  �  	��  �   8�	�A  `e �   >} �K1  r� �
�    �m �
�   $�n �
�   (�m �
�   ,�n �
�   0 qz ��A  8�	`B  `e �   >} �K1  r� �
�    �n �
�   $�m �
�   (;n �
�   ,�n �
�   0 �w ��A  0�	�B  `e �   >} �K1  �n �
�    �m �
�   $��  �
�   ( �x �lB  K   ��B  )top  �G  �  �]  ��B   �	;C  ��  �42   ��  ��B  O{  �
�   ��  �
�   iK  �;C   /  ��  ��B  
AC  ]C  =    	��  �MC  "K   �C  )up  �  �F  �S   FT  
iC  "K   �C  ��   �x  H�  ��  �H   ��  �C  H	�D   `e     >} K1   L� �   %low �  $ +�  �  ( �Z !
�   , r� "
�   0 �f  #�C  4 �f  $�C  8 ��  %�  <%tag &
�   @ *� '�C  D �w )�C  
�D  �D  =    �D  !�  2�D  "K   F�D  �c  +c �c d d �c hc �c  �c P�D  @T	�E   `e V    *� W�D   >} XK1    �}  Y�  ( L� Z�  , ��  ]�   0 �c `�   4 �c c�   8 �y eE  "K   ��E  ��   �s  z�  ��  �T  ܭ   gY  ��E  H�	hF   `e �    *� ��E   >} �K1    �W  ��  ( �}  ��  , L� ��  0 ��  ��  4 ��  �
�   8%tag �
�   < ��  �
�   @  w ��E  
�F  �F  =    hF  !j�  uF  "K   �F  �g  Fe 	h g qf �j �e �f �h i 	�j 
�h ]h  �k 7�F  @E	�G   `e G    *� H�F   ��  I�   >} JK1    ��  K
�   ( }k L
�   , P{  Ml  0 l N�  4 L� O�  8 �x QG  	
  :  	  ;�  �  	��  !M�  	(h  !N�   	l�  !N�   	�  ".�  	�  "/�  	�  "0�  	�  "2�  	w�  "81  	�  "9�  	�  ":�  	�_  ";�   	��  ">�  	�  "J�  	"�  "R�  	t�  "S�   	�w  "T�   	؜  "Y�   	q�  "[�  	Ƚ  "^�  	�  "_�   	�y  "`�   	b�  "c�   	+�  "f�  	��  "i�  	֘ "l�   	�J  "x�   	��  "y�   	ks  "�   	�  "��   	J�  "��   	�i  "��   	��  "��  	��  "��  	��  "��  	<� "��  	��  "��  	��  "��  	5�  "��  	<m  "��   	 K  "��   	�R  "��   	op  "��   	�m  "��   	D  "��   	X�  "��   	If  "��   	� "��   	��  "��  	�U  "��  	`  "��  	J�  "��  	��  "��  	� "�  
L7  CJ  =    	�  "�3J  
�  _J  =    	� "�OJ  
x  {J  =   	 	,�  "�kJ  	R�  "��J  x  
x  �J  =    	�u  "��J  	��  "�q8  	�e  "��   
�   �J  =   � 	(�  "��J  	�  "��  !��  "  !�v  "�   !n�  "�   !4�  "�   !*b "�   !��  "�G  	� #M�   	5 #N�   *�G  '	H_f     +Wz (�   	T_f     *�G  )		P_f     "K   .�K  �y  y  "K   ��K  �x  Qw �v (w �x �w �y �y  ,�x ��K  	@_f     -�/ pMA     �      ��S  .�x �  E 1 .�x �F    .Tw �S  Q M .�v �S  � � .+w �D  � � .�x �S  � � .�w 	�S  9 5 .�y 
�S  s o /3p  �MA      @  �M  0Ap  � � 1@  2Np  � � 3�MA     ur  "M  4Us  5�MA     �u  5�MA     �u  5�MA     �u  5�MA     �u  5�MA     �u  5�MA     �u  5�MA     �u  5�MA     �u  5�MA     �u    /Ho  GNA      �  'HN  0Vo    1�  2co  D B 3LNA     ur  �M  4Us  5QNA     �u  5YNA     �u  5oNA     �u  5wNA     �u  5NA     �u  5�NA     �u  5�NA     �u    /o  �NA      �  0O  0o  k g 1�  2o  � � 3�NA     ur  �N  4Us  5�NA     �u  5�NA     �u  5�NA     �u  5�NA     �u  5�NA     �u  5OA     Mv  5OA     �u  5OA     �u    /�n  HOA      �  9�O  0�n  � � 1�  2�n     3MOA     ur  VO  4Us  5ROA     �u  5hOA     �u  5pOA     �u  5xOA     �u  5�OA     �u  5�OA     �u  5�OA     �u  5�OA     �u  5�OA     �u  5�OA     �u  5�OA     �u    /yn  �OA         F�P  0�n  ) % 1   2�n  a _ 3 PA     ur  9P  4Us  5PA     �u  5PA     �u  5#PA     �u  5+PA     �u  53PA     �u  5;PA     �u    /4n  gPA      `  N+Q  0Bn  � � 1`  2On  � � 3lPA     ur  �P  4Us  5qPA     �u  5�PA     �u  5�PA     �u  5�PA     �u  5�PA     �u  5�PA     �u    /�m  �PA      �  V�Q  0�m  � � 1�  2
n    3�PA     ur  }Q  4Us  5�PA     �u  5�PA     �u  5�PA     �u  5 QA     �u    5vMA     �v  5�MA     ut  3�MA     	y  �Q  4UH4T54Q0 3NA     y  R  4Us  3&NA     !y  R  4Us  50NA     ut  3ANA     	y  NR  4U@4T54Q0 5�NA     ut  3�NA     	y  }R  4U@4T54Q0 51OA     ut  3BOA     	y  �R  4UH4T54Q0 3�OA     y  �R  4Us  3�OA     .y  �R  4Us  5�OA     ut  3�OA     	y  S  4U84T54Q0 5PPA     ut  3aPA     	y  :S  4U84T54Q0 5�PA     ut  3�PA     	y  iS  4U04T54Q0 3QA     y  �S  4Us  6'QA     ;y  4U	��B       �E  �G  �A  `B  �B  -� �KA     d      �X  7th �X  F B 7i ��   � | 8,o  iKA      iKA     >       ��T  0:o  � � 3qKA     qq  MT  4Us  5yKA     �t  5�KA     �t  5�KA     �t  5�KA     �t  5�KA     �t   8�n  �KA      �KA     U       �7U  0�n  � � 3�KA     qq  �T  4Us  5�KA     �t  5�KA     �t  5�KA     �t  5�KA     �t  5�KA     �t  5LA     �u  5LA     �t   8�n  *LA      *LA     l       �V  0�n    32LA     qq  �U  4Us  5FLA     �t  5NLA     �t  5VLA     �t  5^LA     �t  5fLA     �t  5nLA     �t  5vLA     �t  5~LA     �t  5�LA     �t  5�LA     �t   8n  �LA      �LA     A       ��V  0&n  ) ' 3�LA     qq  RV  4Us  5�LA     �t  5�LA     �t  5�LA     �t  5�LA     �t  5�LA     �t   8�m  MA      MA     4       �W  0�m  N L 3MA     qq  �V  4Us  5.MA     �t  56MA     �t  5>MA     �t  5FMA     �t   3dKA     �v  ,W  4U1 5iKA     �s  3�KA     �v  PW  4U2 5�KA     �s  3%LA     �v  tW  4U3 5*LA     �s  5�LA     �v  5�LA     �s  3MA     �v  �W  4U6 5MA     �s  9ZMA     �v  �W  4U7 3aMA     �v  �W  4U0 5fMA     �s  6nMA     qo  4Us     -7. TzHA     �      ��\  .�x V�  y q .Ye WX  � � .�H  XX  & $ .y Y0  M I /Iq  �HA        v?\  0Wq  � � 1  2dq  � � 8�s  �HA      �HA            >�X  5IA     �u   8�s  IA      IA            A,Y  5IA     �u   8�s  +IA      +IA            MaY  50IA     �u   8�s  6IA      6IA            P�Y  5;IA     �u   8�s  AIA      AIA            S�Y  5FIA     �u   8�s  �IA      �IA            q Z  5�IA     �u   8�s  �IA      �IA            �5Z  5�IA     �u   8�s  YJA      YJA     <       ��Z  0�s      5^JA     Mv  5jJA     Mv  5vJA     Mv  5�JA     Mv  5�JA     Mv   8�s  �JA      �JA            ��Z  5�JA     �u   3�HA     ur  �Z  4Us  5�HA     �u  5�HA     �u  5�HA     �u  5IA     �u  5 IA     �u  5(IA     �u  5QIA     �u  5YIA     �u  5aIA     �u  5iIA     �u  5qIA     �u  5yIA     �u  5�IA     �u  5�IA     �u  5�IA     �u  5�IA     �u  5�IA     �u  5�IA     �u  5�IA     �u  5�IA     �u  5�IA     �u  5JA     �u  5JA     �u  5JA     �u  5SJA     �u    5�HA     Gy  5�HA     Sy  5�HA     _y  5�HA     �v  5�HA     ut  3�HA     	y  �\  4U�4T54Q0 3�JA     ky  �\  4Us  3�JA     y  �\  4Us  6KA     ;y  4U	��B       - ( 8�FA     �      �ea  7th :X  8  6  /-q  �FA      �  C-a  0;q  ]  [  8�s  �FA      �FA            ��]  0�s  �  �  5�FA     �t   8�s  �FA      �FA            ��]  0�s  �  �  5�FA     �t   8�s  GA      GA            �^  0�s  �  �  5GA     �t   8�s  GA      GA            �Q^  0�s  �  �  5GA     �t   8�s  GA      GA            ��^  0�s  ! ! 5&GA     �t   8�s  qGA      qGA            ��^  0�s  C! A! 5|GA     �t   8�s  �GA      �GA            �_  0�s  j! h! 5�GA     �t   8�s   HA       HA     <       �_  0�s  �! �! 5,HA     �u  58HA     �u  5DHA     �u  5PHA     �u  5\HA     �u   8�s  \HA      \HA            �_  0�s  �! �! 5gHA     �t   3�FA     qq  �_  4Us  5�FA     �t  5�FA     �t  5�FA     �t  5�FA     �t  5GA     �t  5GA     �t  5.GA     �t  56GA     �t  5>GA     �t  5FGA     �t  5NGA     �t  5VGA     �t  5^GA     �t  5fGA     �t  5qGA     �t  5�GA     �t  5�GA     �t  5�GA     �t  5�GA     �t  5�GA     �t  5�GA     �t  5�GA     �t  5�GA     �t  5HA     �t  5 HA     �t   3�FA     �v  Da  4U1 5�FA     �s  :zHA     �v  4U0  -�) �EA     	      ��b  7i ��   �! �! ;j ��   7sec  K1  v" p" 7li 42  �" �" 7si .2  �" �" 5�EA     Mv  5�EA     Mv  5�EA     Mv  5�EA     Mv  5�EA     Mv  5�EA     Mv  5�EA     Mv  5
FA     Mv  5FA     Mv  5FA     Mv  5?FA     Mv  5IFA     Mv  5TFA     Mv  5]FA     Mv  5fFA     Mv   -�( ��DA     �       ��c  7i ��   # # ;j ��   7sec �K1  �# �# 7li �42  �# �# 7si �.2  $ $ 5�DA     �u  5�DA     �u  5�DA     �u  5�DA     �u  5�DA     �u  5�DA     �u  5�DA     �u  5EA     �u  5EA     �u  5EA     �u  5@EA     �u  5IEA     �u  5REA     �u  5[EA     �u  5dEA     �u   -y' ��AA     �      �ig  7i �
�   <$ :$ /�p  �AA      �  �	[g  <�p  1�  2�p  |$ `$ /�s  �AA      �  �nd  5�AA     �u   8q  BA      BA     C       ��d  <q  5BA     �v  5BA     �v  5&BA     Mv  52BA     Mv  5=BA     �v  5HBA     �v   8�s  �CA      �CA            �e  5�CA     �u   8�s  �CA      �CA            �Se  5�CA     �u   8�p  �CA      �CA     D       �	�e  <�p  =�CA     D       2�p  �% �% 5�CA     �u  5DA     �u  5$DA     �u  5/DA     �u    5BA     �u  5SBA     �u  5^BA     �u  5iBA     �u  5tBA     �u  5BA     �u  5�BA     �u  5�BA     �u  5�BA     �u  5�BA     �u  5�BA     �u  5�BA     �u  5�BA     �u  5�BA     �u  5CA     �u  5CA     �u  54CA     �u  5ICA     �u  5aCA     �u  5lCA     �u  5wCA     �u  5�CA     �u  5�CA     �u  5�CA     �u  5�CA     �u  5�CA     �u  5�CA     �u  5�CA     �u  5�CA     �u  5GDA     �u    5�AA     ut   -" �(?A     �      ��j  7i �
�   �% �% /\p  R?A      �  �	�j  <jp  1�  2wp  & �% /�p  OAA         �	"h  <�p  5sAA     �t  5�AA     �t  5�AA     �t  5�AA     �t   /�s  R?A      P  	Ph  <�s  5_?A     �t   8�p  j?A      j?A     H       �h  <q  5v?A     �v  5�?A     �v  5�?A     �u  5�?A     �u  5�?A     �v  5�?A     �v   8�s  AA      AA            ii  <�s  5AA     �t   8�s  #AA      #AA            r?i  <�s  5.AA     �t   5j?A     �t  5�?A     �t  5�?A     �t  5�?A     �t  5�?A     �t  5�?A     �t  5�?A     �t  5�?A     �t  5@A     �t  5%@A     �t  58@A     �t  5G@A     �t  5Z@A     �t  5e@A     �t  5t@A     �t  5�@A     �t  5�@A     �t  5�@A     �t  5�@A     �t  5�@A     �t  5�@A     �t  5�@A     �t  5�@A     �t  5AA     �t  5AA     �t  5#AA     �t  59AA     �t  5DAA     �t  5OAA     �t  5�AA     �t    5R?A     �s   -$ �?A     
       �k  :(?A     �v  4UM  >�$ �	�  ?A            �Nk  .�| �	�   �& �& 5?A     �v   >�& c	�  ,>A     �       ��l  7i e
�   �& �& 7a f
�  �' �' 7b f�  �' �' 7c f�  �' �' ?Vy g
�l  �@?Qy h
�l  �P5>>A     �v  5T>A     �v  5k>A     wy  3�>A     �y  .l  4Uw 4T@4Q	��B      3�>A     �y  Ll  4Uv 4Tw  5�>A     �v  5�>A     �v  5�>A     �v  5�>A     �v  5�>A     �v  5�>A     �v  5�>A     �v   
�   �l  =    -E CS=A     �       ��m  @�_  C"�   ( ( ?� E
�l  �P7i F	�   k( Y( 5u=A     �v  3�=A     �v  3m  4U0 5�=A     wy  3�=A     �y  jm  4Us 4T@4Q	��B      5�=A     �v  5�=A     �v  5�=A     �v  5�=A     �v  5�=A     �v  5	>A     �v  5>A     �v  5#>A     �v   A�v -�m  Bstr -(�S   A�x n  Bstr '�S  C>} 	�    Ax �4n  Bstr �,�S   A�w �]n  Bstr �+�S  C>} �	�    A~z �yn  Bstr �4�S   Afz ��n  Bstr �3�S  C>} �	�    A>w �n  Bstr (�D   A�w U�n  Bstr U'�D  C>} W	�    A�w 3o  Bstr 32�S   A�x ,o  Bstr 1�S  C>} 	�    A z �Ho  Bstr �,�S   A�y �qo  Bstr �+�S  C>} �	�    Dy �;A     ^       �3p  Estr �.�F  4) .) 3(;A     qq  �o  4Us  50;A     �t  5D;A     �t  5L;A     �t  5T;A     �t  5\;A     �t  5d;A     �t  5l;A     �t  5t;A     �t  F};A     �t   A�v �\p  Bstr �-�F  C>} �	�    A-x �p  Bstr ,?:  ;i 	�    A]y ��p  Bstr �+?:  ;i �	�    Aw g�p  Bstr g,�p   �6  ACz M�p  Bstr M+�p  C�� O	�    A^x 3q  Bstr 3,�G   ABx -q  Bstr +�G   Az �Iq  Bstr �(0   A�z -qq  Bstr -'0  ;pl /	�    D�y ;A            �ur  Estr .X  �) �) /�s  ;A      P   �q  0�s  �) �) 5;A     �t   8�s  ;A      ;A            #r  0�s  �) �) 5;A     �t   Gis  ;A      �  &0vs  "* * G�s  ;A      �  0�s  c* _* F;A     �t     Dx q<A     &       �is  Estr -X  �* �* /�s  q<A      �  �r  5z<A     �u   8�s  <A      <A            s  5�<A     �u   H�s  �<A      �<A            0�s  �* �* I�s  �<A      �<A            �5�<A     �u     J�w ��s  Kstr �.�s   �  J�y ��s  Kstr �-�s   J:y ��s  Kstr �0�J   Jsx ��s  Kstr �/�J   J�w ��s  Kp � R    L.y �R   M�x �};A     +       �ut  Npos �=   /+ -+ OVx �	�   T+ R+ Ni �	�   }+ w+ 5�;A     �y  6�;A     �v  4U0  M�y �H<A     )       ��t  Npos �=   �+ �+ OVx �	�   �+ �+ Ni �	�   , , 5Y<A     �y  5i<A     �v   M�z ��:A     -       ��u  P�| ��   ?, 7, 3�:A     �v  5u  4Us � 3�:A     �v  Pu  4Us 	�$ 3�:A     �v  nu  4U�U@&� :;A     �v  4U�UH%  Q�y ��   <A     7       ��u  O��  �	�   �, �, 5<A     �v  5#<A     �v  5+<A     �v  56<A     �v   M0w z�:A            �Mv  P�| z!l  �, �, 3�:A     �v  ?v  4U�U� F�:A     �v   Q�z pl  �;A            ��v  O��  r	�   :- 4- 5�;A     �v  5<A     �v   J�x c�v  R�| c�   S"y Q�  �v  T��  S
�   U� =�   �<A     �       ��w  P� =�   �- �- V��  ?�   	�e     V5z @1   	 �e     V
w A
�w  �P5=A     �y  3"=A     �y  �w  4Uw 4T 4Q	{�B     4Rs  6F=A     �y  4Q	��B     4Xw   
�   �w  =    U�/ /�   �<A     8       �x  V��  1�   	�e     6�<A     �y  4T	r�B     4Q0  W�v  t:A     R       ��x  0�v  �- �- X�v  �:A            rx  <�v  6�:A     �y  4U	�B       6�:A     �y  4U�l4T14Q1  W�v  �;A     Q       �	y  Y�v  �oZ�;A            �x  [�v  6�;A     �y  4U	5�B       6�;A     �y  4U�o4T14Q1  \� � 
6\3b 3b G]�b �b 	]�t �t <	\��  ��  $7\11 11 q\� � 
7	\Yw Yw F\�d �d �\Q' Q' #K\G�  G�  %/\'�  '�  &\pL pL �\��  ��  'A\[�  [�  f\��  ��  %+^�E �E ( \�L �L �\�K �K � a   �  S#  p{ �*  .QA           k� 9�  �� �  �)  �K   ,	  ^&  �  �1  @�   Q  �    �   	?   62  #	?     &	?   �5  )	?    �@  ,	?   (.  -	?   0*  2�   8;:  5�   < �   1  int �K 8"b   	�  K  �   	�  L  	�  M  
Y   "t  ��  WH  �~  �O  �m  ��   �  ��  ��  	 0t  �  e2    �0  }  ��  t  
Y   J�  D   �C  
D  ���� �C  N�  ڵ  R�  �  	"|  *�  	��  +�  	I�  ,�  	�a  -�  	�  	�   	q  	1  �   t�  
 �   7  
Y   o  �L  M M �L  
Y   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (o  
Y   /�  ��   [r  �4 #�  �   �X  5�  
Y   :b  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K�  
�   P�  =_  ��   R�  N�  ��  ��   �p  Wn  
Y   3�  ��   ({  ��  ğ   F]  8�  
Y   Y  ��   �c  |  ��  l  ��  �   
Y   kj  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {  
Y   ��  &�   �  º  GY  �f  ��   v�  �v  
Y   ��  GQ   ϼ  �  �_  X  &�  �b    	z  ��  "�   E�  #�  e% $�  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�  	� M�   	5 N�   �  =� �  ��  .�  ^�  2s   }�  7y  �� ;Y    	  r�  ,   .� $=  O� )a   &  &  �    �    =  &   2  ?   a  &  Y   `   ?    C  ��  ,�  g  �  oS  '�  dS  ()�  � +
�   � ,&  @�  -
�   >z .
�   �  /`   �H  3�    �   �  K      	�� 7�  	�� 8Y   C  &  K   �'   	��  1&  	]  4C  C  C  Z  K   � I  	Zy  8Z  �  �  K   K   � k  	��  ;�  Ʃ  QY   �  �  �  K     �  	�  W�  �p  #�  �  �   S�  $�  �  �  `    T}  %      `   `    '	K  acv )�  ��  *�  ��  +�   �y -  �Y  6K  ��  :�  s�  <�   �H  =�  xz  >W   c  x @c  
Y   )�  P}  s} z{ �| }} �| d|  | A| �z 	�z 
 9		  x ;
�   y <
�   �{ =�  B		  2�  D
�   ]  E
�  �h  F	�  �N  G	�  �K  H	�  >} J
�   �{ K'	  Q	�	  v1 S
�   v2 T
�  �  U
�  �k V
�  tag W
�  �W  Y
�	  
 �  �	  K    �{ Z�	  �	b
  = �
�   F�  �
�  �~ �	�  h�  �	�  t�  �
�  �k �
�  tag �
�   �| ��	  �	�
  ��  �
�   g{ �
�   �z �n
  �	�
  v1 �
�   v2 �
�  Mp �
�   �  �
�  <p �
�  82  �
�  
 >{ ��
  �	R  x �
�   y �
�  dx �
�  dy �
�  �o �
R  )�  �h   �  h  K   K    �  x  K    %} �   
�	�  x ��   y ��  Mp ��  *� ��  ޽  ��   ~x ��  
Y   (  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  
Y   ��(  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u4  (x	5)   �u z(    � {	�    s |	�    � ~K   N�  �(   ��  �	�    ��  �	�     J]  ��(  5)  S)  K   � !�^  �B)  �   k)  " !�  �`)  #Y   ��,  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  x)  \	.   �Y  	�     *O  	�    ��  	�    �  	�    b�  	�    ��  	�    �  	�    +�  	�    Zp  	�     o�   	�   $ m�  !	�   ( 4�  "	�   , �  #	�   0 �  $	�   4 ��  %	�   8 L� &	�   < ��  '	�   @   (	�   D ��  )	�   H \q *	�   L z�  +	�   P �  ,	�   T /�  -	�   X ʤ  /�,  .  ;.  K   � !��  1+.  �]  ��0  `e ��   x �7  y �7  z �7   ��  �0  (cN  �0  0Mp ��  8�u �(  <� ��   @�H  �0  Hr�  �0  P��  �Y0  X��  �7  `m�  �7  d��  �7  h  �7  l3F  �7  p8F  �7  t=F  �7  x��  ��   |*� ��,  �y� �_0  �s ��   ��� �e0  ��  ��   ��  ��   �ʺ  ��   ��l  ��   �  �  0  � ��  �   � ��  	�   � �R  E2  � f�  �   � I}  �  � ��  0  � H.  Gx  �Y0  >} ��5   �}  ��  �|  ��  
 $0  .  5)  $d  HNE2  mo PV4   ��  QQ;  cmd Rz  �  W7  (_  Y7   #_  [7  $bob ]7  (�  a�   ,�[  b�   0sb  d�   4d]  g];  8�W  hm;  P��  i�  h�� l\4  l�N  mj  |E�  pj  ��W  r};  �~�  s\4  �*� t\4  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �V4  �%�R  ��    %��  ��   %�  ��   %h  ��;  %I�  ��  @ k0  �z H.  	��  ��   	�\  ��  	�  �8   	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  �y  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	,3  x E7   y F7   �{ H3  (T	p3  `e V�   x W7  y X7  z Y7    	�  [83  �a	V4  = c7   F�  d7  �~ e�  h�  f�  
t�  g�  �k h�  tag i�  �N  l
�   ��  oV4  ��  r
\4   iK  up3  0��  x
�   XS�  {V4  `��  ~`   h��  ��   pu| �,5  x K2  �   l4  K    �}  X�,5  v1 ��5   v2 ��5  dx �7  dy �7  �  ��  �k ��  tag ��  �W  ��	  �o ��5  $��  ��5  4SX  ��5  8d�  ��5  @��  �
�   H��  �`   P 25  l4  �z �|3  �	�5  2�  �7   ]  �7  �h  ��  �N  ��  
�K  ��  >} ��5   85  �}  �D5  
Y   ��5  ��   �  o�  ��   ��  ��5  ,3  7  �5  K    �u  �l4  �z �$0  8�	6  v1 ��5   v2 ��5  82  �7  Mp ��  [�  �6   �  ��6   SX  ��5  (d�  ��5  0 �5  �5  A{ �6  4	�6  &x 7   &y 	7  &dx 
7  &dy 7   �o �6   )�  h  0 7  7  K   K    (} �6  �  *�  'v  @2�7   @�  4�7   &x1 5�   &x2 6�    .]  87   5]  97   �� :7   ��  =�    �  @7    ��  C7  $ �n  G�7  ( 9x  H�7  0 �^  I�7  8 �6  �  >�  K 7  '�h  PR�8   s�  U�8    �H  V�8  &x1 X�   &x2 Y�   &gx \7  &gy ]7  &gz `7   &gzt a7  $ �x  d7  ( � f7  , ~�  i7  0 t  k7  4 .� l�   8 �  p�8  @ 	�  r�   H �7  7  �h  t�7  �	9   �c  ��    �O  �9   �x  �
(9   �  (9  K    �  89  K    I�  ��8  �	l9   �  ��     �  �l9   89  �  �E9  (��	):     �7    �  �	�    t�  �	�    ��  �	�    /�  �	�    �  �	�  &top �	):  )��  �	�  U)��  �	�  V)� �	):  W)�  �	�  � �  ::  K   ? ��  �9  	�:  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %G:  �:  �:  K    	S�  '�:  
Y   7�:  {�   U�  ~�   >	$;  �� @e0   s A
�   sx B7  sy C7   Nz E�:  
Y   1Q;  ��   ��  ��   �y  90;  �   m;  K    �  };  K    �  �;  K    $;  �;  K    hy �k0  (�	<  in ��   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
\4  �a  �
�   $ ��  ��;  ��	�<  2�  �
�    I�  ��  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��<  ( <  �<  K    ޴  �<  	.L  &�<  7  	׮  )�<  	�  +�<  	�  ,�<  	�Q  .�8  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7L=  �   	��  8L=  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�=  r9  	��  H�   	��  I�5  	��  K�   	a� L�7  	w�  N�   	P{ O�5  	��  Q�   	��  R >  6  	��  T�   	�� U>  7  	�}  W�   	u| X�6  	M�  Z�   	P�  [6  	��  a7  	��  b7  	�  c7  	�p  e�  	�T  f�>  �;  	�a  j�  �   �>  K   � 	ը  l�>  �  �>  K   @ 	�p  m�>  	 �  p7  	p|  q�  	$Y  v�   	�K  y�   	g  {?  ::  	d�  |?  	��   7  		�  !7  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +7  	`�  ,7  	A�  -7  	��  /�   	��  1�   	P�  2�   �8  �?  K   K   / 	��  E�?  �8  �?  K   / 	Ԁ  F�?  �8  @  K   K    	7� G�?  	�R  I�   	��  J�8  	��  U�   	P�  \�  	��  ]�  	L�  ^�  	ߵ  _�  	�  a�  	@�  �7  	[�  6  	 �  �6  	SX  �5  	d�  �5  	��  �   	_�   �   	��  "�  	��  %�  	'�  &�  	�]  (�  �7  A  K   � 	�P  *�@  	ӯ  +&A  �7  	|  -8A  �8  	��  .8A  	��  /8A  \A  lA  �   �    	��  �7  �   VA  	qY  "xA  	�  #xA  �  �A  K   ? 	��  %�A  	��  &�A  7  �A  K   � 	@Y  (�A  7  �A  K   ? 	V�  )�A  �8  B  K    	�h   �A  	�   &B  �8  	�   �8  	�f   !�A  	r�   "�A  	��   %�7  	��   &�7  	׆   '7  	��   (7  	�   *7  	��   +7  	�  !�8  	��  !�   	�_  !�   	�_  !�   	b  !7  	t  !7  	j�  !"y  	�  !:�   	��  !;�   	��  !<�   	�W  !>�8  	hn  !@7  	U~  !A7  	�  !B7  	 �  !C7  	%�  !Fy  	�u  !Hy  	z  !Iy  	ʓ  "C�  �  �C  K    	��  "b|C  �   �C  K    	��  "c�C  	0K  "d�   	?�  "e�   "�	D  x "�7   y "�7  dx "�7  dy "�7   ��  "��C  "�2D  �p "�
V4  ��  "�
�6   "�	aD  {q "�7   ��  "��  d "�	D   t�  "�2D  aD  }D  K   � 	r "�mD  	�T  "��D  aD  	l�  "�7  	�  "�7  	?k  "�7  	�d  "�7  	2~ "�D  	��  "��  	��  "�7  	k�  "�7  	Z�  "��6  �6  E  K    	�v  "�E  	�v  "��   	"�  "�V4  !�  "y  !�U  "�7  !��  "�7  !t�  "�   !�  "	�   !.Y  "
7  !7Y  "7  !�h  "�E  V4  !*� "\4  !<i  "\4  	G  #�  	��  #�   �   �E  K    
Y   #�F  *top  �G  �  �]  #��E   #�	cF  ��  #��6   ��  #�F  O{  #�
�   ��  #�
�   iK  #�cF   p3  ��  #�F  iF  �F  K    	��  #�uF  #Y   #�F  *up  �  �F  �S   FT  #
�F  #Y   #�F  ��   �x  H�  ��  �H   ��  #�F  H#	�G   `e #�    >} #�5   L� #7   &low #7  $ +� # 7  ( �Z #!
�   , r� #"
�   0 �f  ##�F  4 �f  #$�F  8 ��  #%�  <&tag #&
�   @ *� #'�F  D �w #) G  �G  �G  K    �G  !�  #2�G  #Y   #�H  ��   �s  z�  ��  �T  ܭ   gY  #��G  H#�	�H   `e #��    *� #�H   >} #��5    �W  #�7  ( �}  #�7  , L� #�7  0 ��  #��  4 ��  #�
�   8&tag #�
�   < ��  #�
�   @  w #�$H  �H  �H  K    �H  !j�  #�H  ) $�H  J @$�I  � $"�    � $'
�E  �� $*	�   
 $-�I  �9 $0	�    Ml  $3	�   $	
 $8	�   (C� $;	�   ,� $?	�   0� $B`   8 �H   $H	�I  � $K�    C� $N	�   "8 $Q`   t $T`    . $V�I  	: $��   	3 $��   	� $��   	� $��   	O $��   	�
 $��   �H  *J  " 	R %J  �I  AJ  " 	� %6J  	 &V�   z  	��  'M�  	(h  'N�   	l�  'N�   	�  (.�  	�  (/�  	�  (0�  	�  (2�  	w�  (8�  	�  (9�  	�  (:b  	�_  (;�   	��  (>�  	�  (J�  	"�  (R�  	t�  (S�   	�w  (T�   	؜  (Y�   	q�  ([�  	Ƚ  (^�  	�  (_�   	�y  (`�   	b�  (c�   	+�  (f�  	��  (i�  	֘ (l�   	�J  (x�   	��  (y�   	ks  (�   	�  (��   	J�  (��   	�i  (��   	��  (��  	��  (��  	��  (��  	<� (��  	��  (��  	��  (��  	5�  (��  	<m  (��   	 K  (��   	�R  (��   	op  (��   	�m  (��   	D  (��   	X�  (��   	If  (��   	� (��   	��  (��  	�U  (��  	`  (��  	J�  (��  	��  (��  	� (��  �;  �L  K    	�  (��L  �  M  K    	� (��L  �  #M  K   	 	,�  (�M  	R�  (�;M  �  �  QM  K    	�u  (�AM  	��  (��<  	�e  (��   �   �M  K   � 	(�  (�uM  	�  (��  !��  (�  !�v  (�   !n�  (�   !4�  (�   !*b (�   !��  (YJ  +�=  3	h_f     +�=  4	�_f     +�=  6	�`f     +�=  7		x`f     +�=  9	p`f     +�=  :	``f     +�=  <	�_f     +�=  =	`_f     +>  ?	@`f     +>  @
	X`f     +$>  B	0`f     +0>  C
	8`f     +<>  E	h`f     +H>  F
	�_f     ,p| H�   	��e     +bE  R	l`f     +oE  S	�`f     +UE  T		P`f     +HE  V		�_f     +|E  X
	H`f     +�E  Y
	D`f     +�E  [
	�`f     +;E  e	�`f     +#M  k	�_f     +/M  l	(`f     +QM  m	 `f     -� O#^A            �P  .)^A     �_  ..^A     �_  /9^A     `   -8! �\[A     �      ��S  0K% ��   ". . 1map ��   �. �. 0�| ��   �. �. 0  ��   / �. 2i �
�   =/ 9/ 3� �
�E  ��4C� �
�   {/ u/ 5�S  �\A     �\A     �       '@R  6�S  �/ �/ 7�\A     �       8�S  �/ �/ 8�S  '0 %0 9�S  ]A         �	�Q  6T  L0 J0 6	T  s0 o0 :   8#T  �0 �0 8.T  /1 '1 8;T  �1 �1 8HT  2 �1 ;UT  �@<{]A     `  �Q  =T	�B     =Qs =R@ >�]A     `  =U	V�B        <�\A     )`  �Q  =U|  <�\A     5`  R  =U| =T5 <�\A     A`  *R  =T5=Q	�`f      >]A     M`  =U|    .�[A     Y`  <�[A     e`  iR  =U5=T6 .�[A     q`  <(\A     }`  �R  =U��=T9 <Q\A     �`  �R  =U�� <e\A     �U  �R  =Uv
 <q\A     �^  �R  =Uv <y\A     [  �R  =Uv <�\A     �V  S  =Uv <�\A     �W  %S  =Uv <�\A     (\  =S  =Uv <�\A     �Y  US  =Uv <�\A     ]  mS  =Uv .�\A     sT  <�]A     �X  �S  =Uv <�]A     �`  �S  =Us  .
^A     �`  .^A     �`   ?�} ��S  @C� ��   A/} �	�   A	| �	�    ?{| �cT  @s �"y  Blen �6Y   Ci �Y   A[| �Y   A`5 �y  A�| �Y   A-| �cT   Y   sT  K    -�| !YA     ?      ��U  4�| #�U  ?2 =2 2i $�   z2 b2 2j %�   y3 u3 2li &�6  �3 �3 4>} '�5  4 �3 2ss ( >  �4 z4 2seg )�7  �4 �4 3�o *�5  �@4�� +�   55 %5 <�YA     A`  `U  =T5=Q0 <sZA     �`  xU  =Uw  <�ZA     �`  �U  =Uw  >�ZA     �`  =Uw   �6  -L| ��XA     �       ��V  0�O  ��   6 6 Di �	�    4r� �	�   e6 a6 4	| �	�   �6 �6 <�XA     )`  -V  =Us  <�XA     A`  IV  =T5=Q0 <�XA     M`  aV  =Us  >YA     A`  =Us =T5=Q0  -!{ ��WA     �       ��W  0�O  ��   �6 �6 4"8 �y  -7 +7 2i ��   X7 P7 2msd ��W  �7 �7 2sd �6  '8 !8 <�WA     )`  W  =Uv  <�WA     A`  :W  =T5=Q}  < XA     5`  WW  =Uv =T1 <;XA     �`  oW  =Us  <JXA     �`  �W  =Us <]XA     �`  �W  =Usr E�XA     �`  =U�U  	  -X{ �VA     �      ��X  0�O  ��   z8 r8 4"8 �y  �8 �8 2i ��    9 �8 2mld ��X  '9 #9 2ld ��6  _9 ]9 2v1 ��5  �9 �9 2v2 ��5  �9 �9 <)VA     )`  �X  =U|  <JVA     A`  �X  =T5=Q}  <sVA     5`  �X  =U| =T1 .�VA     �`  E�WA     �`  =U�U  �	  - | OjUA     �       ��Y  0�O  O�   �9 �9 4"8 Qy  ": : 2i R�   ^: X: 2mt S;M  �: �: 3	} T�  �F47| U�   �: �: 4_t V�  6; 4; <�UA     5`  �Y  =Uv =T1 <�UA     )`  �Y  =Uv  <�UA     �`  �Y  =U�F >VA     �`  =Uv   -g} *�TA     �       � [  0�O  *�   b; Z; 4"8 ,y  �; �; 2i -
�   �; �; 2j .
�   '< !< 2k /
�   w< s< 2mn 0 [  �< �< 2no 1>  �< �< <�TA     )`  �Z  =Us  <�TA     A`  �Z  =T5=Q0 <�TA     5`  �Z  =Us =T1 EjUA     �`  =U�U  x  -Y} 	�SA     �       �"\  0�O  	�   = �< 4"8 y  b= `= 2i �   �= �= 2ms "\  �= �= 2ss �5  \> V> <�SA     )`  �[  =U|  <�SA     A`  �[  =T5=Q}  <"TA     5`  �[  =U| =T1 <YTA     a  �[  =Us  <jTA     a  \  =Usn E�TA     �`  =U�U  b
  FG{ �8SA     �       �]  G�O  ��   �> �> H"8 �y  ? ? Ii ��   Q? I? Ims �]  �? �? Iss � >  D@ :@ <@SA     )`  �\  =Us  <\SA     A`  �\  =T5=Q0 <oSA     5`  �\  =Us =T1 E�SA     �`  =U�U  �
  F�z ��QA     C      �N^  G�O  ��   �@ �@ H"8 �y  <A :A Ii ��   aA _A Iml �N^  �A �A Ili ��7  �A �A H�| ��6  �A �A H �  ��   JB HB J<p ��   H�W  ��   {B wB <RA     )`  �]  =Uv  <'RA     A`  ^  =T5=Q}  <ORA     5`  +^  =Uv =T1 .SA     T^  E8SA     �`  =U�U  �
  K�| ��5  �^  ,�{ ��  	��e     ,9} �85  	 �e      F| v.QA     p       �w_  G�O  v�   �B �B H"8 xy  C C Ii y�   EC =C Iml zw_  �C �C Ili {�5  GD =D <6QA     )`  (_  =Us  <UQA     A`  D_  =T5=Q0 <hQA     5`  a_  =Us =T1 E�QA     �`  =U�U  	  LT^  �QA     W       ��_  :�  <�QA     a  �_  =U0=T	 �e     =Q4 >�QA     a  =U4=T	$�e     =Q4   M{ { #�M�| �| #'	M0{ 0{  6MF�  F�  bM� � 	!M�} �} ?M� � BM� � 6M{ { @	M�| �| &/ME} E} 8	MYw Yw "FM[�  [�  fM�{ �{ =M�% �% M�} �} #*	M�{ �{ )%M�L �L &M�L �L )Mw! w! )0M} } I	MH_  H_  
#	M�s �s ,M) ) )+M�H �H *;	 �G   ��  S#  �} �*  9^A     #      �� J�  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �  
K   Y�  ��   �c  |  ��  l  ��  �   
K   k   _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {�  
K   �_  &�   �  º  GY  �f  ��   v�  �,  
K   ��  GQ   ϼ  �  �_  X  &�  �b    	0  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�  B  t�  	 �   C  O  e  =   �' T  	��  
1e  	]  
4�  O  O  �  =   � �  	Zy  
8�  �  �  =   =   � �  	��  
;�  Ʃ  
QK   �  �  �  =     �  	�  
W�  �p  #       S�  $)  /  :  R    T}  %F  L  \  R   R    '	�  acv )  ��  *  ��  +:   �y -\  �Y  6�  ��  :�  s�  <�   �H  =�  xz  >�   �  x @�  B  �  =    4  	  =    
�	P  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x �	  
K   �  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �\  
K   �@"  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�  (x	�"  �u z�   � {	�   s |	�   � ~�  N�  @"  ��  �	�   ��  �	�     J]  �M"  �"  �"  =   � �^  ��"  �   �"    �  ��"  !K   �I&  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �"  \	�'  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /V&  �'  �'  =   � ��  1�'  �]  ���)  `e ��   x �C  y �C  z �C   ��  ��)  (cN  ��)  0Mp ��  8�u ��  <� ��   @�H  ��)  Hr�  ��)  P��  ��)  X��  �C  `m�  �C  d��  �C  h  �C  l3F  �C  p8F  �C  t=F  �C  x��  ��   |*� �I&  �y� ��)  �s ��   ��� ��)  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  �)  ���  �   ���  	�   ��R  �+  �f�  �   �I}  P  ���  �)  � �'  Gx  ��)  >} �./   �}  �B  �|  �B  
 �)  �'  �"  "d  HN�+  mo P�-   ��  Q�4  cmd R0  �  WC  (_  YC   #_  [C  $bob ]C  (�  a�   ,�[  b�   0sb  d�   4d]  g�4  8�W  h�4  P��  iy  h�� l�-  l�N  m   |E�  p   ��W  r5  �~�  s�-  �*� t�-  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��-  �#�R  ��    #��  ��   #�  ��   #h  �5  #I�  �y  @ �)  �z �'  �  	��  ��   	�\  �y  	�  �,  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  ��+  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	�,  x EC   y FC   �{ H�,  (T	-  `e V�   x WC  y XC  z YC    	�  [�,  �a	�-  = cC   F�  dC  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  o�-  ��  r
�-   iK  u-  0��  x
�   XS�  {�-  `��  ~R   h��  ��   pu| ��.  x �+  �   �-  =    �}  X��.  v1 �s/   v2 �s/  dx �C  dy �C  �  �B  �k �B  tag �B  �W  ��  �o �y/  $��  �g/  4SX  �./  8d�  �./  @��  �
�   H��  �R   P �.  �-  �z �-  �	./  2�  �C   ]  �C  �h  �B  �N  �B  
�K  �B  >} �./   �.  �}  ��.  
K   �g/  ��   �  o�  ��   ��  �@/  �,  C  �/  =    �u  ��-  �z ��)  8�	0  v1 �s/   v2 �s/  82  �C  Mp ��  [�  �0   �  �0   SX  �./  (d�  �./  0 4/  �/  A{ ��/  4	�0  $x C   $y 	C  $dx 
C  $dy C  �o �0  )�  �  0 C  �0  =   =    (} )0  �  *�  %v  @2g1  @�  4g1   $x1 5�   $x2 6�   .]  8C  5]  9C  �� :C  ��  =�   �  @C   ��  CC  $�n  Gm1  (9x  Hm1  0�^  Im1  8 0  B  >�  K�0  %�h  PR\2  s�  U\2   �H  V\2  $x1 X�   $x2 Y�   $gx \C  $gy ]C  $gz `C   $gzt aC  $�x  dC  (� fC  ,~�  iC  0t  kC  4.� l�   8�  pb2  @	�  r�   H �1  �0  �h  t�1  �	�2  �c  �y   �O  ��2  �x  �
�2   B  �2  =    �  �2  =    I�  �u2  �	�2  �  ��    �  ��2   �2  �  ��2  &��	�3    �C   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  $top �	�3  '��  �	�  U'��  �	�  V'� �	�3  W'�  �	�  � �  �3  =   ? ��  �3  	14  ~�  _   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�3  14  M4  =    	S�  '=4  
K   7z4  {�   U�  ~�   >	�4  �� @�)   s A
�   sx BC  sy CC   Nz Ez4  
K   1�4  ��   ��  ��   �y  9�4  �   �4  =    y  5  =    y  5  =    �4  /5  =    hy ��)  	.L  &G5  C  	׮  )G5  	�  +G5  	�  ,G5  	�Q  .b2  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�5  �   	��  8�5  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F6  3  	��  H�   	��  Is/  	��  K�   	a� Lg1  	w�  N�   	P{ O./  	��  Q�   	��  Rm6  �/  	��  T�   	�� U�6  �0  	�}  W�   	u| X0  	M�  Z�   	P�  [0  	��  aC  	��  bC  	�  cC  	�p  e�  	�T  f�6  /5  	�a  j�  �    7  =   � 	ը  l7  �  =7  =   @ 	�p  m,7  	 �  pC  	p|  q�  	$Y  v�   	�K  y�   	g  {�7  �3  	d�  |�7  	��   C  		�  !C  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +C  	`�  ,C  	A�  -C  	��  /�   	��  1�   	P�  2�   b2  =8  =   =   / 	��  E'8  b2  Y8  =   / 	Ԁ  FI8  b2  {8  =   =    	7� Ge8  	�R  I�   	��  Jb2  	��  U�   	P�  \<  	��  ]<  	L�  ^<  	ߵ  _<  	�  a<  	@�  g1  	[�  0  	 �  0  	SX  ./  	d�  ./  	��  �   	_�   �   	��  "y  	��  %y  	'�  &y  	�]  (y  s1  {9  =   � 	�P  *k9  	ӯ  +�9  s1  	|  -�9  b2  	��  .�9  	��  /�9  �9  �9  �   �    	��  m1  �   �9  	qY  "�9  	�  #�9  B  :  =   ? 	��  %	:  	��  &	:  C  B:  =   � 	@Y  (2:  C  _:  =   ? 	V�  )N:  h2  {:  =    	�h  k:  	�  �:  h2  	�  h2  	�f  !	:  	r�  "	:  	��  %m1  	��  &m1  	׆  'C  	��  (C  	�  *C  	��  +C  	�  b2  	��  �   	�_  �   	�_  �   	b  C  	t  C  	j�  "�+  	�  :�   	��  ;�   	��  <�   	�W  >b2  	hn  @C  	U~  AC  	�  BC  	 �  CC  	%�  F�+  	�u  H�+  	z  I�+  	ʓ  C�  P  �;  =    	��  b�;  �   <  =    	��  c<  	0K  d�   	?�  e�   �	q<  x �C   y �C  dx �C  dy �C   ��  �9<  ��<  �p �
�-  ��  �
0   �	�<  {q �C   ��  �y  d �	}<   t�  ��<  �<  �<  =   � 	r ��<  	�T  �=  �<  	l�  �C  	�  �C  	?k  �C  	�d  �C  	2~ �q<  	��  �y  	��  �C  	k�  �C  	Z�  �0  0  �=  =    	�v  �t=  	�v  ��   	"�  ��-  �  �+  �U  m1  ��  m1  t�  �   �  	�   .Y  
C  7Y  C  �h  >  �-  *� �-  <i  �-  	G  y  	��  �   
K   �i>  (top  �G  �  �]  �H>   �	�>  ��  �0   ��  �i>  O{  �
�   ��  �
�   iK  ��>   -  ��  �u>  �>  �>  =    	��  ��>  !K   ?  (up  �  �F  �S   FT  
�>  !K   P?  ��   �x  H�  ��  �H   ��  "?  H	@  `e �   >} ./  L� C   $low C  $+�  C  (�Z !
�   ,r� "
�   0�f  #?  4�f  $?  8��  %y  <$tag &
�   @*� 'P?  D �w )]?  -@  -@  =    @  �  2@  !K   �t@  ��   �s  z�  ��  �T  ܭ   gY  �@@  H�	A  `e ��   *� �t@  >} �./   �W  �C  (�}  �C  ,L� �C  0��  �y  4��  �
�   8$tag �
�   <��  �
�   @  w ��@  5A  5A  =    A  j�  %A  )�}  
C  	�`f     )�o !
C  	�`f     )�q "
C  	�`f     )1~ $q<  	�`f     *t2x %
C  	�`f     *t2y &
C  	�`f     �   �A  =    )�} (�A  	�`f     +�f -y  �aA     �       ��B  ,t1 .�-  �D �D ,t2 /�-  .E (E -s1 1
�   ~E zE -s2 2
�   �E �E .F� 3
�   �E �E .�} 4
�   8F 2F .~ 5
�   �F �F /SbA     �B   +"~ 	y  �`A     �       �[C  0~ �   �F �F -bsp �6  lG fG .<p 
�   �G �G /�`A     [C  1+aA     gF  9C  2Qs  3AaA     �B  4YaA     gF  2Qq   5�} �	y  _A     �      ��E  6num ��   #H H 7seg �g1  qH oH 8��  �0  �H �H 7s1 ��   �H �H 7s2 ��   bI \I 8r� ��   �I �I 7sub �m6  �I �I 8g� �./  �I �I 8� �./  J J 8l�  �C  AJ ?J 8�  �C  fJ dJ 9�} �q<  ��7v1 �s/  �J �J 7v2 �s/  �J �J 8{q �C  �J �J 8�  �C  (K $K 1=_A     �G  �D  2U	j�B     2Ts  1�_A     gF  �D  2U| 2Tv 2Qq  1�_A     gF  "E  2U{ 2Tz 2Qq  1�_A     gF  :E  2Qq  1`A     gF  RE  2Qq  1h`A     �E  xE  2U	�`f     2T�� 1�`A     �G  �E  2T��� 3�`A     �G   5~ fC  �^A     s       �aF  6v2 gaF  hK ^K 6v1 haF  �K �K 9{q jC  V7num kC  `L \L 7den lC  �L �L 3�^A     �G  3�^A     �G  3�^A     �G  3�^A     �G  /
_A     �G   q<  :�} 0�   �F  ;x 1C  ;y 2C  <=� 3aF  =dx 5C  =dy 6C  >Ϸ  7C  >�T  8C   ?gF  9^A     h       ��G  @xF  M M @�F  EM AM A�F  QB�F  �M ~M B�F  �M �M B�F  #N !N B�F  HN FN CgF  P  @�F  mN kN @�F  �N �N @xF  �N �N DP  E�F  E�F  E�F  E�F     F��  ��  7FH_  H_  	#	Fd  d  	"	 Pb   t�  S#  �~ �*  \bA           �� ��  �)  �=   ,	  int ^&  9�  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2D   8;:  5D   < �   1  �K 8"b   	�  K
  �   	�  L
  	�  M
  0t  4  e2    �0  }  ��  (  
[   J�  D   �C  
D  ���� �C  N\  ڵ  RP  �  
[   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
[   /!  ��   [r  �4 #�  �   �X  5�  
[   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K-  
D   P�  =_  ��   R�  N�  ��  ��   �p  W�  
[   3  ��   ({  ��  ğ   F]  8�  
[   YG  ��   �c  |  ��  l  ��  �   
[   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {G  
[   ��  &�   �  º  GY  �f  ��   v�  ��  
[   �  GQ   ϼ  �  �_  X  &�  �b   �   ,  =    I  <  =    ;  L  =    
	�	�  x 	�I   y 	�I  Mp 	�I  *� 	�I  ޽  	�I   ~x 	�L  
 	+  ��  
"B   E�  
#B  e% 
$I  u  
%
�  �8 
&
�  ��  
)
�  /b  
-
�  ��  
.	D   a  
2
�  �T  
3
�   Mx 
4�  �  D   =  +  	��  M�  	(h  ND   	l�  ND   	�  ~�  �   �S  
D   ��   
D     !
D   �g  "
D   �^  #
D    ��  %t  �  �  =    	S�  '�  t�   D   �       =   �'   	��  1  	]  43        J  =   � 9  	Zy  8J  �  q  =   =   � [  	��  ;q  Ʃ  Q[   �  �  �  =     �  	�  W�  �p  #D  S�  $�  �  �  K    T}  %�  �     K   K    '	.  acv )�  ��  *�  ��  +�   �y -   �Y  6.  ��  :{  s�  <{   �H  ={  xz  >:   F  x @F  
[   �
  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  
[   �q$  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�
  (x	�$  �u z�
   � {	D   s |	D   � ~.  N�  q$  ��  �	D   ��  �	D     J]  �~$  �$  	%  =   � �^  ��$  �   !%    �  �%  ![   �z(  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  .%  \	�)  �Y  	D    *O  	D   ��  	D   �  	D   b�  	D   ��  	D   �  	D   +�  	D   Zp  	D    o�   	D   $m�  !	D   (4�  "	D   ,�  #	D   0�  $	D   4��  %	D   8L� &	D   <��  '	D   @  (	D   D��  )	D   H\q *	D   Lz�  +	D   P�  ,	D   T/�  -	D   X ʤ  /�(  �)  �)  =   � ��  1�)  
[   7*  {�   U�  ~�   >	[*  �� @[*   s A
D   sx B�  sy C�   �$  Nz E*  �]  ��C,  `e ��   x ��  y ��  z ��   ��  �C,  (cN  �C,  0Mp ��  8�u ��
  <� �D   @�H  �C,  Hr�  �C,  P��  �~,  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  �D   |*� �z(  �y� ��,  �s �D   ��� �[*  ��  �D   ��  �D   �ʺ  �D   ��l  �D   � �  C,  ���  D   ���  	D   ��R  d.  �f�  D   �I}  �  ���  C,  � m*  Gx  �~,  >} ��8   �}  �I  �|  �I  
 I,  �)  "d  HNd.  mo P�.   ��  Q�.  cmd R+  �  W�  (_  Y�   #_  [�  $bob ]�  (�  aD   ,�[  bD   0sb  dD   4d]  g�.  8�W  h�.  P��  i�  h�� l�.  l�N  m�  |E�  p�  ��W  r�.  �~�  s�.  �*� t�.  ��� wD   ���  xD   �X�  |D   ��e  D   ���  �D   �g  �D   ��u  �D   �|G ��   �Q  �D   ��  �D   �o�  ��.  �#�R  �D    #��  �D   #�  �D   #h  �/  #I�  ��  @ �,  �z m*  
[   1�.  ��   ��  ��   �y  9w.  
[   @�.  el �l �l  j.  D   �.  =    �  �.  =    D   �.  =    �  /  =    a*  /  =    hy ��,  (�	�/  in ��   d  �
D   �x  �
D   D  �
D   5O  �
D   �� �
�.  �a  �
D   $ ��  �'/  ��	00  2�  �
D    I�  ��  r�  �
D   �H  �
D   *F  �
D   ��  �
D   	�  �
D   ѵ  �
D   ��  �
D    F� �
D   $�  �00  ( �/  @0  =    ޴  ��/  	�  .�  	�  /�  	�  0�  	�  2�  	w�  8!  	�  9�  	�  :�  	�_  ;�   	��  >�  	�  J�  	"�  R�  	t�  SD   	�w  TD   	؜  YD   	q�  [�  	Ƚ  ^�  	�  _D   	�y  `D   	b�  cD   	+�  f�  	��  i�  	֘ lD   	�J  xD   	��  yD   	ks  D   	�  �D   	J�  �D   	�i  �D   	��  ��  	��  ��  	��  ��  	<� ��  	��  ��  	��  ��  	5�  ��  	<m  �D   	 K  �D   	�R  �D   	op  �D   	�m  �D   	D  �D   	X�  �D   	If  �D   	� �D   	��  ��  	�U  ��  	`  ��  	J�  ��  	��  ��  	� �  /  �2  =    	�  ��2  �  �2  =    	� ��2  �  �2  =   	 	,�  ��2  	R�  �3  �  �  3  =    	�u  �
3  	��  �@0  	�e  ��   �   O3  =   � 	(�  �>3  	�  ��  ��    �v  D   n�  D   4�  D   *b D   ��  J  	"|  *�  	��  +�  	I�  ,�  	�a  -�  �3  $
[   "14  ��  WH  �~  �O  �m  ��   �  ��  ��  	 	�  D   	q  I4  �   =� [4  ��  .�4  ^�  25   }�  77  �� ;[    	�4  r�  �4   .� $�4  O� )5   %�4  �4  �    O4  �4  �4  �4   �4  %1   5  �4  [   K   1    �4  ��  ,�4  5  oS  '/5  dS  ()�5  � +
   � ,�4  @�  -
D   >z .
D   �  /K   �H  3�5    #5  	�� 7�5  	�� 8[   	��  ��   	�\  ��  	�  ��5  �  	��  �D   	��  �D   	2�  ��  	��  �D   	Ɇ  �7  	��  �D   	��  �D   	�h  �D   	rK  �D   	l�  �D   	]�  �D   	��  �D   C	�6  x E�   y F�   �{ Hd6  (T	�6  `e V�   x W�  y X�  z Y�    	�  [�6  �a	�7  = c�   F�  d�  �~ eI  h�  fI  
t�  gI  �k hI  tag iI  �N  l
D   ��  o�.  ��  r
�.   iK  u�6  0��  x
D   XS�  {�.  `��  ~K   h��  �D   pu| �n8  x �}  X�n8  v1 �#9   v2 �#9  dx ��  dy ��  �  �I  �k �I  tag �I  �W  �,  �o �)9  $��  �9  4SX  ��8  8d�  ��8  @��  �
D   H��  �K   P t8  �7  �z ��6  �	�8  2�  ��   ]  ��  �h  �I  �N  �I  
�K  �I  >} ��8   z8  �}  ��8  
[   �9  ��   �  o�  ��   ��  ��8  �6  �  99  =    �u  ��7  �z �I,  8�	�9  v1 �#9   v2 �#9  82  ��  Mp ��  [�  ��9   �  ��9   SX  ��8  (d�  ��8  0 �8  99  A{ �Q9  4	2:  &x �   &y 	�  &dx 
�  &dy �  �o 2:  )�  <  0 �  H:  =   =    (} �9  �  *�  'v  @2;  @�  4;   &x1 5D   &x2 6D   .]  8�  5]  9�  �� :�  ��  =D   �  @�   ��  C�  $�n  G;  (9x  H;  0�^  I;  8 �9  I  >�  Kb:  '�h  PR<  s�  U<   �H  V<  &x1 XD   &x2 YD   &gx \�  &gy ]�  &gz `�   &gzt a�  $�x  d�  (� f�  ,~�  i�  0t  k�  4.� lD   8�  p<  @	�  rD   H 0;  U:  �h  t0;  �	Z<  �c  ��   �O  �Z<  �x  �
j<   I  j<  =    �  z<  =    I�  �%<  �	�<  �  �D    �  ��<   z<  �  ��<  (��	k=    ��   �  �	D   t�  �	D   ��  �	D   /�  �	D   �  �	�  &top �	k=  )��  �	�  U)��  �	�  V)� �	k=  W)�  �	�  � �  |=  =   ? ��  ��<  	.L  &�=  �  	׮  )�=  	�  +�=  	�  ,�=  	�Q  .<  	��  0D   	��  1D   	(_  2D   	դ  4D   	�j  7>  D   	��  8>  	@�  <D   	�O  =D   	(g  >D   	�^  ED   	�u FU>  �<  	��  HD   	��  I#9  	��  KD   	a� L;  	w�  ND   	P{ O�8  	��  QD   	��  R�>  E9  	��  TD   	�� U�>  H:  	�}  WD   	u| X�9  	M�  ZD   	P�  [�9  	��  a�  	��  b�  	�  c�  	�p  e�  	�T  fK?  /  	�a  j�  D   n?  =   � 	ը  l]?  �  �?  =   @ 	�p  mz?  	 �  p�  	p|  q�  	$Y  vD   	�K  yD   	g  {�?  |=  	d�  |�?  	��   �  		�  !�  	�3 #D   	_  $D   	-�  (D   	�f  )D   	�G  +�  	`�  ,�  	A�  -�  	��  /D   	��  1D   	P�  2D   <  �@  =   =   / 	��  Eu@  <  �@  =   / 	Ԁ  F�@  <  �@  =   =    	7� G�@  	�R  ID   	��  J<  	��  UD   	P�  \�3  	��  ]�3  	L�  ^�3  	ߵ  _�3  	�  a�3  	@�  ;  	[�  �9  	 �  �9  	SX  �8  	d�  �8  	��  D   	_�   D   	��  "�  	��  %�  	'�  &�  	�]  (�  #;  �A  =   � 	�P  *�A  	ӯ  +�A  #;  	|  -�A  <  	��  .�A  	��  /�A  B  'B  D   D    	��  ;  �   B  	qY  "3B  	�  #3B  I  hB  =   ? 	��  %WB  	��  &WB  �  �B  =   � 	@Y  (�B  �  �B  =   ? 	V�  )�B  <  �B  =    	�h   �B  	�   �B  <  	�   <  	�f   !WB  	r�   "WB  	��   %;  	��   &;  	׆   '�  	��   (�  	�   *�  	��   +�  	�  !<  	��  !D   	�_  !D   	�_  !D   	b  !�  	t  !�  	j�  !"7  	�  !:D   	��  !;D   	��  !<D   	�W  !><  	hn  !@�  	U~  !A�  	�  !B�  	 �  !C�  	%�  !F7  	�u  !H7  	z  !I7  	ʓ  "C�  �  GD  =    	��  "b7D  D   cD  =    	��  "cSD  	0K  "dD   	?�  "eD   "�	�D  x "��   y "��  dx "��  dy "��   ��  "��D  "��D  �p "�
�.  ��  "�
�9   "�	E  {q "��   ��  "��  d "�	�D   t�  "��D  E  8E  =   � 	r "�(E  	�T  "�PE  E  	l�  "��  	�  "��  	?k  "��  	�d  "��  	2~ "��D  	��  "��  	��  "��  	k�  "��  	Z�  "��9  �9  �E  =    	�v  "��E  	�v  "�D   	"�  "��.  �  "7  �U  ";  ��  ";  t�  "D   �  "	D   .Y  "
�  7Y  "�  �h  "^F  �.  *� "�.  <i  "�.  	G  #�  	��  #D   �   �F  =    
[   #��F  *top  �G  �  �]  #��F   #�	G  ��  #��9   ��  #��F  O{  #�
D   ��  #�
D   iK  #�G   �6  ��  #��F  $G  @G  =    	��  #�0G  ![   #sG  *up  �  �F  �S   FT  #
LG  ![   #�G  ��   �x  H�  ��  �H   ��  #�G  H#	nH  `e #�   >} #�8  L� #�   &low #�  $+� # �  (�Z #!
D   ,r� #"
D   0�f  ##sG  4�f  #$sG  8��  #%�  <&tag #&
D   @*� #'�G  D �w #)�G  �H  �H  =    nH  �  #2{H  ![   #F�H  �c  +c �c d d �c hc �c  ![   #�I  ��   �s  z�  ��  �T  ܭ   gY  #��H  H#�	�I  `e #��   *� #�I  >} #��8   �W  #��  (�}  #��  ,L� #��  0��  #��  4��  #�
D   8&tag #�
D   <��  #�
D   @  w #�I  �I  �I  =    �I  j�  #�I  ![   #DJ  �g  Fe 	h g qf �j �e �f �h i 	�j 
�h ]h  �k #7�I  ![   #=mJ  1l  �k  @#E	�J  `e #G�   *� #HDJ  ��  #I�  >} #J�8   ��  #K
D   (}k #L
D   ,P{  #MI  0l #N�  4L� #O�  8 �x #QmJ  	� $MD   	5 $ND   ) %'K  J @%�K  � %"�    � %'
�F  �� %*	D   
 %-�K  �9 %0	D    Ml  %3	D   $	
 %8	D   (C� %;	D   ,� %?	D   0� %BK   8 K   %H	�K  � %K�    C� %N	D   "8 %QK   t %TK    . %V�K  	: %�D   	3 %�D   	� %�D   	� %�D   	O %�D   	�
 %��   K  ZL    	R &OL  �K  qL    	� &fL  
[   &r O  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	 'VD   7	wO  �~ 9�   �  :
D   8~ ;
D   �~ <
D   L� =
D    �~ ?,O  D	�O  �~ F
D    I G
�F  �~ H
�F  L� I
D    � J�O  wO  �O  =    	�� P�O  	� Q�O  wO  �O  P  =    + `�O  	�[e     ,�O  �		 af     ,�O  �
	�`f     	� �I  �9  _P  =   ? 	& �OP  -~F  B
	�cf     -�F  C	�`f     .CP  Y	�`f     ._P  Z
	�cf     /�} ^�mA     �      ��Q  0>} `�8  �N �N 1i a
D   O �N 2:nA     �`  Q  3Us  2OnA     �`  ,Q  3Us  2`nA     �`  NQ  3Us 3T?3Q0 2pnA     �`  fQ  3Us  2�nA     �`  ~Q  3Us  2�nA     �`  �Q  3Us 3Tv  2�nA     �`  �Q  3Us  4�nA     �`  3U	��B       5~~ �D   �kA     $      ��T  6��  ��9  �O �O 1s1 ��8  'P %P 1s2 ��8  RP JP 1s3 ��8  �P �P 0�k �D   Q �P 1rtn �D   iQ cQ 1i �D   �Q �Q 0�v ��T  �Q �Q 0: ��  VR RR 0�~ �I  �R �R 7�T  VlA     VlA     �       '�S  8�T  �R �R 8�T  �R �R 8�T  S S 8�T  FS DS 9VlA     �       :OU  ;\U  clA     �       <]U  rS nS 2�lA     a  vS  3U	��B     3T2 2�lA     a  �S  3T	��e      2�lA     a  �S  3T	��e      4�lA     a  3T	�B     3RF    2�kA     gZ  �S  3Uu 3T|  2�kA     x^  T  3Uu 3Ts  2lA     +a  2T  3U	*�B      2VlA     +a  QT  3U	��B      2$mA     6a  sT  3U@3T63Q0 2/mA     Ba  �T  3Uv  2pmA     6a  �T  3U@3T63Q0 4{mA     Ba  3Uv   �J  =� �jU  >: �#�=  >�~ �:;  >��  �"�9  > �2�8  ?�~ �D   	�[e     ?6 �D   	��e     ?�~ �D   	��e     � �D   @Ap �D     /�~ E?jA     _      �V  0� G�O  �S �S 1pic H
D   �S �S 1i I
D   T �S 0��  J�9  �T �T BYjA     Na  4kA     Za  3Us3TG  /Q �eiA     �       ��V  6�R  �)K?  U U 0>} ��8  �U �U C�iA     fa  B�iA     sa  2$jA     fa  �V  3T03Q03RD C0jA     Na  D=jA     �`  3U	��B       /�o ��hA     k       �~W  6�p ��.  �V �V 6��  ��9  ?W 3W 1ok �
D   �W �W 23iA     a  )W  3Us 3T3 2BiA     �a  FW  3Us 3T3 2XiA     �a  hW  3Us 3T33Q0 DciA     �a  3U�T  /�q ��eA     F      ��Y  6� �D   �W �W 6<p �D   ;Y 'X 6�p ��.  �d Xd 0��  ��9  zi Ti 1ok �
D   �j �j 2YfA     �a  X  3Us  2�fA     �a  5X  3Us  2�fA     �a  MX  3Us  2gA     �a  jX  3Us 3T1 CgA     Na  2*gA     �a  �X  3Us  2AgA     �a  �X  3Us  2\gA     �a  �X  3Us  2gA     �a  �X  3Us  2�gA     �a  �X  3Us  C�gA     
b  2�gA     b  Y  3Us  2�gA     a  ,Y  3Us  2�gA     �a  DY  3Us  C�gA     �a  ChA     �a  ChA     �a  C/hA     �a  CphA     �a  C�hA     �a  C�hA     b  C�hA     a   5�m �D   ~eA     6       �gZ  6>} ��8  !k k Emax �D   �k }k 1i �
D   �k �k 1min �
D   %l !l 0��  ��9  ]l [l 0Wy ��8  �l �l 4�eA     x^  3Uu 3Tx   5Vb �D   JeA     4       ��Z  F��  ��9  U6' �D   �l �l 1i �	D   m m  5nb �	�  eA     5       �g[  Esec �3�8  Zm Rm 1i �
D   �m �m 0Wy ��9  n n 0�  ��8  Ln Jn 0  ��  sn on 45eA     x^  3Uu 3Tx   5Ic ��  �dA     8       �\  Esec �*�8  �n �n 1i �D   o o 0Wy ��9  wo uo 0�  ��8  �o �o 0  ��  �o �o 4 eA     x^  3Uu 3Tx   5�k J�  DdA     �       �]  Esec K�8  p p 6� LD   �p �p 1i ND   q �p 1h OD   �q �q 1min PD   r r 0Wy Q�9  7r 5r 0�  R�8  fr br 0  S�  �r �r ? T]  ��~2udA     x^  ]  3Uu 3T}  4�dA     �`  3U	��B       �  .]  =    5Nk (	�  dA     7       ��]  Esec (1�8  �r �r 1i *D   Bs :s 0Wy +�9  �s �s 0�  ,�8  �s �s 0�v -�  �s �s 40dA     x^  3Uu 3Tx   5l 	�  �cA     4       �x^  Esec 0�8  :t 2t 1i D   �t �t 0Wy �9  �t �t 0�  �8  ,u *u 0�v �  Qu Ou 4�cA     x^  3Uu 3Tx   G�m ��8  �cA            ��^  H��  ��9  UIsec ��8  T Gtk �D   �cA     !       ��^  J>} �D   xu tu H��  �D   T G�k ��8  pcA     2       �O_  J� �D   �u �u H��  �D   TH<p �D   Q Glk ��9  BcA     .       ��_  J� �D   �u �u H��  �D   TH<p �D   Q K�| �\bA     �       ��`  Li �
D   9~bA     �       M�~ ��   1v +v MI ��   |v zv 2�bA     #b  `  3Uv  2�bA     /b  3`  3U|  2�bA     /b  K`  3Uv  B�bA     ;b  2�bA     Gb  p`  3U|  2�bA     Gb  �`  3Uv  4cA     �`  3U	��B     3Tv 3Q|    Nlm lm #�	N�m �m #�NJn Jn #�	O"d "d #}	O�c �c #�N(n (n #�	N��  ��  (7N��  ��  %NSJ SJ )"	NF�  F�  bP�E �E , N� � 6N3b 3b "GN�. �. $<N� � '6Odj dj "N� � *!OUf Uf #nO�c �c #rO�t �t #7Ni i #�Nmn mn #�	N^n ^n #�O@b @b #O�t �t #>	O�b �b #N�n �n #�	O�k �k #iN�# �# $=O�~ �~ #xNe~ e~ +1Nw! w! +0Nj j <N) ) ++ �R   �  S#  f� �*  joA           � Ŕ  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �   	"  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�  4  	"|  *y  	��  +y  	I�  ,y  	�a  -y  
K   	�  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  	(e  
K   	/�  ��   [r  �4 #�  �   �X  	5�  
K   	:X  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  	K�  
�   	P�  =_  ��   R�  N�  ��  ��   �p  	Wd  
K   
3�  ��   ({  ��  ğ   F]  
8�  
K   
Y  ��   �c  |  ��  l  ��  �   
K   
k`  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  
{  
K   
��  &�   �  º  GY  �f  ��   v�  
�l  
K   
��  GQ   ϼ  �  �_  X  &�  �b   t�   �   �  �    =   �' �  	��  1  	]  4#  �  �  :  =   � )  	Zy  8:  �  a  =   =   � K  	��  ;a  Ʃ  QK   r  ~  �  =     �  	�  W�  �p  #�  �  �   S�  $�  �  �  R    T}  %�  �  �  R   R    '	+  acv )�  ��  *�  ��  +�   �y -�  �Y  6+  ��  :x  s�  <x   �H  =x  xz  >7   C  x @C  B  �  =    4  �  =    
�	�  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x ��  
K   N
  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  
K   ��#  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  uZ
  (x	[$  �u zN
   � {	�   s |	�   � ~+  N�  �#  ��  �	�   ��  �	�     J]  ��#  [$  y$  =   �  �^  �h$  �   �$  !  �  ��$  "K   ��'  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �$  \	D)  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /�'  D)  a)  =   �  ��  1Q)  �]  ��D+  `e �~   x ��  y ��  z ��   ��  �D+  (cN  �D+  0Mp �r  8�u �N
  <� ��   @�H  �D+  Hr�  �D+  P��  �+  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� ��'  �y� ��+  �s ��   ��� ��+  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  D+  ���  �   ���  	�   ��R  k-  �f�  �   �I}  �  ���  D+  � n)  Gx  �+  >} ��0   �}  �B  �|  �B  
 J+  D)  [$  #d  HNk-  mo P�/   ��  Q�6  cmd R"  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g�6  8�W  h�6  P��  iy  h�� l�/  l�N  m`  |E�  p`  ��W  r�6  �~�  s�/  �*� t�/  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��/  �$�R  ��    $��  ��   $�  ��   $h  ��6  $I�  �y  @ �+  �z n)  �  	��  ��   	�\  �y  	�  ��-  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  �~-  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	_.  x E�   y F�   �{ H?.  (T	�.  `e V~   x W�  y X�  z Y�    	�  [k.  �a	�/  = c�   F�  d�  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  o�/  ��  r
�/   iK  u�.  0��  x
�   XS�  {�/  `��  ~R   h��  ��   pu| �_0  x q-  �   �/  =    �}  X�_0  v1 �1   v2 �1  dx ��  dy ��  �  �B  �k �B  tag �B  �W  ��  �o �1  $��  �1  4SX  ��0  8d�  ��0  @��  �
�   H��  �R   P e0  �/  �z ��.  �	�0  2�  ��   ]  ��  �h  �B  �N  �B  
�K  �B  >} ��0   k0  �}  �w0  
K   �1  ��   �  o�  ��   ��  ��0  _.  �  *1  =    �u  ��/  �z �J+  8�	�1  v1 �1   v2 �1  82  ��  Mp �r  [�  ��1   �  ��1   SX  ��0  (d�  ��0  0 �0  *1  A{ �B1  4	#2  %x �   %y 	�  %dx 
�  %dy �  �o #2  )�  �  0 �  92  =   =    (} �1  �  *�  &v  @23  @�  43   %x1 5�   %x2 6�   .]  8�  5]  9�  �� :�  ��  =�   �  @�   ��  C�  $�n  G3  (9x  H3  0�^  I3  8 �1  B  >�  KS2  &�h  PR�3  s�  U�3   �H  V�3  %x1 X�   %x2 Y�   %gx \�  %gy ]�  %gz `�   %gzt a�  $�x  d�  (� f�  ,~�  i�  0t  k�  4.� l�   8�  p4  @	�  r�   H !3  F2  �h  t!3  �	K4  �c  �y   �O  �K4  �x  �
[4   B  [4  =    �  k4  =    I�  �4  �	�4  �  ��    �  ��4   k4  �  �x4  '��	\5    ��   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  %top �	\5  (��  �	�  U(��  �	�  V(� �	\5  W(�  �	�  � �  m5  =   ? ��  ��4  	�5  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %z5  �5  �5  =    	S�  '�5  
K   76  {�   U�  ~�   >	W6  �� @�+   s A
�   sx B�  sy C�   Nz E6  
K   1�6  ��   ��  ��   �y  9c6  �   �6  =    y  �6  =    y  �6  =    W6  �6  =    hy ��+  (�	@7  in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�/  �a  �
�   $ ��  ��6  ��	�7  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��7  ( @7  �7  =    ޴  �L7  	.L  &8  �  	׮  )8  	�  +8  	�  ,8  	�Q  .4  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  78  �   	��  88  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�8  �4  	��  H�   	��  I1  	��  K�   	a� L3  	w�  N�   	P{ O�0  	��  Q�   	��  R39  61  	��  T�   	�� UQ9  92  	�}  W�   	u| X�1  	M�  Z�   	P�  [�1  	��  a�  	��  b�  	�  c�  	�p  er  	�T  f�9  �6  	�a  jr  �   �9  =   � 	ը  l�9  r  :  =   @ 	�p  m�9  	 �  p�  	p|  qr  	$Y  v�   	�K  y�   	g  {K:  m5  	d�  |K:  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   4  ;  =   =   / 	��  E�:  4  ;  =   / 	Ԁ  F;  4  A;  =   =    	7� G+;  	�R  I�   	��  J4  	��  U�   	P�  \.  	��  ].  	L�  ^.  	ߵ  _.  	�  a.  	@�  3  	[�  �1  	 �  �1  	SX  �0  	d�  �0  	��  �   	_�   �   	��  "y  	��  %y  	'�  &y  	�]  (y  3  A<  =   � 	�P  *1<  	ӯ  +Y<  3  	|  -k<  4  	��  .k<  	��  /k<  �<  �<  �   �    	��  3  �   �<  	qY  "�<  	�  #�<  B  �<  =   ? 	��  %�<  	��  &�<  �  =  =   � 	@Y  (�<  �  %=  =   ? 	V�  )=  	4  A=  =    	�h  1=  	�  Y=  	4  	�  	4  	�f  !�<  	r�  "�<  	��  %3  	��  &3  	׆  '�  	��  (�  	�  *�  	��  +�  	�  4  	��  �   	�_  �   	�_  �   	b  �  	t  �  	j�  "~-  	�  :�   	��  ;�   	��  <�   	�W  >4  	hn  @�  	U~  A�  	�  B�  	 �  C�  	%�  F~-  	�u  H~-  	z  I~-  	ʓ  C~  �  �>  =    	��  b�>  �   �>  =    	��  c�>  	0K  d�   	?�  e�   �	7?  x ��   y ��  dx ��  dy ��   ��  ��>  �e?  �p �
�/  ��  �
�1   �	�?  {q ��   ��  �y  d �	C?   t�  �e?  �?  �?  =   � 	r ��?  	�T  ��?  �?  	l�  ��  	�  ��  	?k  ��  	�d  ��  	2~ �7?  	��  �y  	��  ��  	k�  ��  	Z�  ��1  �1  J@  =    	�v  �:@  	�v  ��   	"�  ��/   �  ~-   �U  3   ��  3   t�  �    �  	�    .Y  
�   7Y  �   �h  �@  �/   *� �/   <i  �/  	G  y  	��  �   �	?A  F� �
?A   L� �
?A  	K% �B   �   OA  =    -� �A  
K   �|A  )top  �G  �  �]  �[A   �	�A  ��  ��1   ��  �|A  O{  �
�   ��  �
�   iK  ��A   �.  ��  ��A  �A  �A  =    	��  ��A  "K   (B  )up  �  �F  �S   FT  
B  "K   cB  ��   �x  H�  ��  �H   ��  5B  H	#C  `e ~   >} �0  L� �   %low �  $+�  �  (�Z !
�   ,r� "
�   0�f  #(B  4�f  $(B  8��  %y  <%tag &
�   @*� 'cB  D �w )pB  @C  @C  =    #C   �  20C  "K   F�C  �c  +c �c d d �c hc �c  "K   ��C  ��   �s  z�  ��  �T  ܭ   gY  ��C  H�	kD  `e �~   *� ��C  >} ��0   �W  ��  (�}  ��  ,L� ��  0��  �y  4��  �
�   8%tag �
�   <��  �
�   @  w ��C  �D  �D  =    kD   j�  xD  "K   �D  �g  Fe 	h g qf �j �e �f �h i 	�j 
�h ]h  "K   =E  1l  �k  	� M�   	5 N�   ) 9E  J @�E  � "�    � '
?A  �� *	�   
 -�E  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 -E   H	F  � K�    C� N	�   "8 QR   t TR    . V�E  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   -E  lF  ! 	R  aF  F  �F  ! 	�  xF  
K    r2I  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	 !V�   "  	��  "My  	(h  "N�   	l�  "N�   	�  #.y  	�  #/y  	�  #0y  	�  #2y  	w�  #8�  	�  #9�  	�  #:X  	�_  #;�   	��  #>y  	�  #Jy  	"�  #R�  	t�  #S�   	�w  #T�   	؜  #Y�   	q�  #[y  	Ƚ  #^�  	�  #_�   	�y  #`�   	b�  #c�   	+�  #fy  	��  #iy  	֘ #l�   	�J  #x�   	��  #y�   	ks  #�   	�  #��   	J�  #��   	�i  #��   	��  #�y  	��  #�y  	��  #�y  	<� #�y  	��  #�y  	��  #�y  	5�  #�y  	<m  #��   	 K  #��   	�R  #��   	op  #��   	�m  #��   	D  #��   	X�  #��   	If  #��   	� #��   	��  #�y  	�U  #�y  	`  #�y  	J�  #�y  	��  #�y  	� #��  �6  �K  =    	�  #��K  y  �K  =    	� #��K  �  L  =   	 	,�  #��K  	R�  #� L  �  �  6L  =    	�u  #�&L  	��  #��7  	�e  #��   �   kL  =   � 	(�  #�ZL  	�  #�y   ��  #�   �v  #�    n�  #�    4�  #�    *b #�    ��  #>I  OA  �L  =   ( *q� *�L  	`^e     �   M  =   c *[� ]�L  	�gf     *:� ^�   	�gf     +�A  _	�ef     ,�i y  �qA     �      �uO  -�p �/  w �v -��  �1  +{ #{ -<p �   �{ �{ .JrA     �Q  �M  /Us /T�U .YrA     �Q  �M  /Us  .prA      R  �M  /Us  .|rA     uO  N  /Us /T0 0�rA     R  .�rA     R  7N  /Us  .�rA     %R  ON  /Us  .�rA     2R  gN  /Us  .�rA     uO  �N  /Us /T0 0 sA     ?R  .9sA     KR  �N  /Us  .ksA     XR  �N  /Us /T6 .�sA     KR  �N  /Us  .�sA     2R  �N  /Us /T0 .-tA     R  O  /Us  .?tA     %R  +O  /Us  .QtA     XR  HO  /Us /T6 .jtA     eR  `O  /Us  1wtA     uO  /Us   2i �{pA     Z      �ZP  3��  ��1  �{ �{ 3R� �	�   e| [| 4�� ��   �| �| 4� ��   /} )} 4� ��   ~} x} 5i ��   �} �} 4*u ��   �~ �~ 0�pA     qR  08qA     qR  0�qA     qR  6�qA     ZP  /U�U  7� ��P  8��  ��1  9w �|A  8P{  ��   8{� ��   :i �
�    2{ ejoA     �       �%Q  5i g
�   �~ �~ 4�8 h
�     4K% i
�   � � .�oA     }R  Q  /Uv  1�oA     }R  /Uv	  ;ZP  �oA     ~       ��Q  <gP  � � <sP  W� Q� <}P  �� �� <�P  �� �� =�P  I� G� >ZP   pA     Z       ?�P  ?}P  ?sP  ?gP  @ pA     Z       =�P  s� m� 6zpA     �R  /U	(�B         A�c �c mA�k �k iB~~ ~~ rB�. �. <A�t �t 7AUf Uf nA@b @b B�# �# =A�c �c rA7d 7d wB^n ^n �B� � !6Bw! w! $0B��  ��  %7 �M   ��  S#  �� �*  �tA     �      � ��  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �  
K   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
K   /  ��   [r  �4 #�  �   �X  5�  
K   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K&  
�   P�  =_  ��   R�  N�  ��  ��   �p  W�  
K   3�  ��   ({  ��  ğ   F]  8�  
K   kX  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {  
K   ��  &�   �  º  GY  �f  ��   v�  �d  B  �  =    4  �  =    
	�	
  x 	�B   y 	�B  Mp 	�B  *� 	�B  ޽  	�B   ~x 	��  
 	�  ��  
";   E�  
#;  e% 
$B  u  
%
�  �8 
&
�  ��  
)
�  /b  
-
�  ��  
.	�   a  
2
�  �T  
3
�   Mx 
4  �  �   �  �  	��  My  	(h  N�   	l�  N�   	C  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�  C  _  =    	S�  'O  t�   �   k  w  �  =   �' |  	��  1�  	]  4�  w  w  �  =   � �  	Zy  8�  �  �  =   =   � �  	��  ;�  Ʃ  QK   �      =     
  	�  W  �p  #�  S�  $D  J  U  R    T}  %a  g  w  R   R    '	�  acv ),  ��  *8  ��  +U   �y -w  �Y  6�  ��  :�  s�  <�   �H  =�  xz  >�   �  x @�  
K   U
  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �  
K   ��#  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  ua
  (x	b$  �u zU
   � {	�   s |	�   � ~�  N�  �#  ��  �	�   ��  �	�     J]  ��#  b$  �$  =   � �^  �o$  �   �$    �  ��$  !K   ��'  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �$  \	K)  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /�'  K)  h)  =   � ��  1X)  >	�)  �� @�)   s A
�   sx Bk  sy Ck   b$  Nz Eu)  
K   p�*  �! 9& +! v( %# 0  B& @�! ��"  w#  	$  �-  S%  �)   0  @&  ��"    !0    m0    b-    �.    �$     /   @ %   � <"    U-    5'    	!  �]  ��y,  `e ��   x �k  y �k  z �k   ��  �y,  (cN  �y,  0Mp ��  8�u �U
  <� ��   @�H  �y,  Hr�  �y,  P��  ��,  X��  �k  `m�  �k  d��  �k  h  �k  l3F  �k  p8F  �k  t=F  �k  x��  ��   |*� ��'  �y� ��,  �s ��   ��� ��)  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  y,  ���  �   ���  	�   ��R  �.  �f�  �   �I}  
  ���  y,  � �*  Gx  ��,  >} �';   �}  �B  �|  �B  
 ,  K)  "d  HN�.  mo P�.   ��  Q�.  cmd R�  �  Wk  (_  Yk   #_  [k  $bob ]k  (�  a�   ,�[  b�   0sb  d�   4d]  g�.  8�W  h�.  P��  iy  h�� l /  l�N  mX  |E�  pX  ��W  r/  �~�  s /  �*� t /  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��.  �#�R  ��    #��  ��   #�  ��   #h  � /  #I�  �y  @ �,  �z �*  
K   1�.  ��   ��  ��   �y  9�.  �.  �   �.  =    y   /  =    �   /  =    y   /  =    �)  0/  =    hy ��,  (�	�/  in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
 /  �a  �
�   $ ��  �</  ��	E0  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  �E0  ( �/  U0  =    ޴  ��/  	�  .y  	�  /y  	�  0y  	�  2y  	w�  8  	�  9�  	�  :�  	�_  ;�   	��  >y  	�  Jy  	"�  R�  	t�  S�   	�w  T�   	؜  Y�   	q�  [y  	Ƚ  ^�  	�  _�   	�y  `�   	b�  c�   	+�  fy  	��  iy  	֘ l�   	�J  x�   	��  y�   	ks  �   	�  ��   	J�  ��   	�i  ��   	��  �y  	��  �y  	��  �y  	<� �y  	��  �y  	��  �y  	5�  �y  	<m  ��   	 K  ��   	�R  ��   	op  ��   	�m  ��   	D  ��   	X�  ��   	If  ��   	� ��   	��  �y  	�U  �y  	`  �y  	J�  �y  	��  �y  	� ��  0/  �2  =    	�  ��2  y  �2  =    	� ��2  
  3  =   	 	,�  ��2  	R�  �3  
  
  /3  =    	�u  �3  	��  �U0  	�e  ��   �   d3  =   � 	(�  �S3  	�  �y  ��  �  �v  �   n�  �   4�  �   *b �   ��  �  ) �3  J @f4  � "�    � '
f4  �� *	�   
 -v4  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 �   v4  =    �3   H	�4  � K�    C� N	�   "8 QR   t TR    . V|4  $�4  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��   �3   5    	R 5  �4  75    	� ,5  
K   r�7  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	 V�   	��  ��   	�\  �y  	�  �8  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  ��  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	�8  x Ek   y Fk   �{ H�8  (T	9  `e V�   x Wk  y Xk  z Yk    	�  [�8  �a	�9  = ck   F�  dk  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  o�.  ��  r
 /   iK  u9  0��  x
�   XS�  {�.  `��  ~R   h��  ��   pu| ��:  x �}  X��:  v1 �l;   v2 �l;  dx �k  dy �k  �  �B  �k �B  tag �B  �W  ��  �o �r;  $��  �`;  4SX  �';  8d�  �';  @��  �
�   H��  �R   P �:  �9  �z �9  �	';  2�  �k   ]  �k  �h  �B  �N  �B  
�K  �B  >} �';   �:  �}  ��:  
K   �`;  ��   �  o�  ��   ��  �9;  �8  k  �;  =    �u  ��9  �z �,  8�	
<  v1 �l;   v2 �l;  82  �k  Mp ��  [�  �
<   �  �<   SX  �';  (d�  �';  0 -;  �;  A{ ��;  4	{<  %x k   %y 	k  %dx 
k  %dy k  �o {<  )�  �  0 k  �<  =   =    (} "<  �  *�  &v  @2`=  @�  4`=   %x1 5�   %x2 6�   .]  8k  5]  9k  �� :k  ��  =�   �  @k   ��  Ck  $�n  Gf=  (9x  Hf=  0�^  If=  8 <  B  >�  K�<  &�h  PRU>  s�  UU>   �H  VU>  %x1 X�   %x2 Y�   %gx \k  %gy ]k  %gz `k   %gzt ak  $�x  dk  (� fk  ,~�  ik  0t  kk  4.� l�   8�  p[>  @	�  r�   H y=  �<  �h  ty=  �	�>  �c  �y   �O  ��>  �x  �
�>   B  �>  =    �  �>  =    I�  �n>  �	�>  �  ��    �  ��>   �>  �  ��>  '��	�?    �k   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  %top �	�?  (��  �	�  U(��  �	�  V(� �	�?  W(�  �	�  � �  �?  =   ? ��  �
?  	.L  &�?  k  	׮  )�?  	�  +�?  	�  ,�?  	�Q  .[>  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7P@  �   	��  8P@  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�@  �>  	��  H�   	��  Il;  	��  K�   	a� L`=  	w�  N�   	P{ O';  	��  Q�   	��  RA  �;  	��  T�   	�� U"A  �<  	�}  W�   	u| X<  	M�  Z�   	P�  [
<  	��  ak  	��  bk  	�  ck  	�p  e�  	�T  f�A  0/  	�a  j�  �   �A  =   � 	ը  l�A  �  �A  =   @ 	�p  m�A  	 �  pk  	p|  q�  	$Y  v�   	�K  y�   	g  {B  �?  	d�  |B  	��   k  		�  !k  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +k  	`�  ,k  	A�  -k  	��  /�   	��  1�   	P�  2�   [>  �B  =   =   / 	��  E�B  [>  �B  =   / 	Ԁ  F�B  [>  C  =   =    	7� G�B  	�R  I�   	��  J[>  	��  U�   	P�  \�4  	��  ]�4  	L�  ^�4  	ߵ  _�4  	�  a�4  	@�  `=  	[�  
<  	 �  <  	SX  ';  	d�  ';  	��  �   	_�   �   	��  "y  	��  %y  	'�  &y  	�]  (y  l=  D  =   � 	�P  *D  	ӯ  +*D  l=  	|  -<D  [>  	��  .<D  	��  /<D  `D  pD  �   �    	��  f=  �   ZD  	qY  "|D  	�  #|D  B  �D  =   ? 	��  %�D  	��  &�D  k  �D  =   � 	@Y  (�D  k  �D  =   ? 	V�  )�D  a>  E  =    	�h  E  	�  *E  a>  	�  a>  	�f  !�D  	r�  "�D  	��  %f=  	��  &f=  	׆  'k  	��  (k  	�  *k  	��  +k  	�  [>  	��  �   	�_  �   	�_  �   	b  k  	t  k  	j�  "�  	�  :�   	��  ;�   	��  <�   	�W  >[>  	hn  @k  	U~  Ak  	�  Bk  	 �  Ck  	%�  F�  	�u  H�  	z  I�  	ʓ   C�  
  �F  =    	��   b�F  �   �F  =    	��   c�F  	0K   d�   	?�   e�    �	G  x  �k   y  �k  dx  �k  dy  �k   ��   ��F   �6G  �p  �
�.  ��   �
<    �	eG  {q  �k   ��   �y  d  �	G   t�   �6G  eG  �G  =   � 	r  �qG  	�T   ��G  eG  	l�   �k  	�   �k  	?k   �k  	�d   �k  	2~  �G  	��   �y  	��   �k  	k�   �k  	Z�   �<  <  H  =    	�v   �H  	�v   ��   	"�   ��.  �   �  �U   f=  ��   f=  t�   �   �   	�   .Y   
k  7Y   k  �h   �H  �.  *�   /  <i    /  	G  !y  	��  !�   
K   !� I  )top  �G  �  �]  !��H   !�	WI  ��  !�<   ��  !� I  O{  !�
�   ��  !�
�   iK  !�WI   9  ��  !�I  ]I  yI  =    	��  !�iI  !K   !�I  )up  �  �F  �S   FT  !
�I  !K   !�I  ��   �x  H�  ��  �H   ��  !�I  H!	�J  `e !�   >} !';  L� !k   %low !k  $+� ! k  (�Z !!
�   ,r� !"
�   0�f  !#�I  4�f  !$�I  8��  !%y  <%tag !&
�   @*� !'�I  D �w !)�I  �J  �J  =    �J  �  !2�J  !K   !�K  ��   �s  z�  ��  �T  ܭ   gY  !��J  H!�	�K  `e !��   *� !�K  >} !�';   �W  !�k  (�}  !�k  ,L� !�k  0��  !�y  4��  !�
�   8%tag !�
�   <��  !�
�   @  w !�K  �K  �K  =    �K  j�  !�K  *�~ *�   �tA     �      ��M  +��  +<  ā �� +<p ,�   �� �� +�p -�.  .� "� ,i /
�   Ƃ �� ,tag 0
�   y� s� ,m 1�.  ރ ڃ ,fog 2�.  � � ,an 3K   P� N� -`e 4�M  u� s� ->} 5';  �� �� -�p 6k  Ą �� -�p 7k  �� �� -�� 8k  8� 4� ..uA     �M  M  /Us  .puA     �M  BM  /U| /T} /Q~ /R' .}uA     �M  ZM  /T# .�uA     �M  rM  /R' 0�uA     �M  /T#  �  1;i ;i  �	1�( �(  k1� � 6 )I   W�  S#  ŀ �*  vA     �       $ �  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �  t�   �   �  �  �  =   �' �  	��  1�  	]  4�  �  �  �  =   � �  	Zy  8�  �    =   =   � �  	��  ;  Ʃ  QK   $  0  F  =     5  	�  WF  
K   	�  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  	(W  
K   	/�  ��   [r  �4 #�  �   �X  	5�  
K   	:J  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  	K�  
�   	P�  =_  ��   R�  N�  ��  ��   �p  	WV  
K   
3�  ��   ({  ��  ğ   F]  
8�  
K   
Y  ��   �c  |  ��  l  ��  �   
K   
kR  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  
{  
K   
��  &�   �  º  GY  �f  ��   v�  
�^  
K   
��  GQ   ϼ  �  �_  X  &�  �b   �p  #�  �  �   S�  $�      R    T}  %    .  R   R    '	\  acv )�  ��  *�  ��  +   �y -.  �Y  6\  ��  :�  s�  <�   �H  =�  xz  >h   t  x @t  B  �  =    4  �  =    
�	"  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x ��  
K   	  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �.  
K   �#  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�	  (x	�#  �u z	   � {	�   s |	�   � ~\  N�  #  ��  �	�   ��  �	�     J]  �#  �#  �#  =   � �^  ��#  �   �#    �  ��#  !K   �'  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �#  \	u(  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /('  u(  �(  =   � ��  1�(  �]  ��u*  `e ��   x ��  y ��  z ��   ��  �u*  (cN  �u*  0Mp �$  8�u �	  <� ��   @�H  �u*  Hr�  �u*  P��  ��*  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� �'  �y� ��*  �s ��   ��� ��*  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  u*  ���  �   ���  	�   ��R  �,  �f�  �   �I}  "  ���  u*  � �(  Gx  ��*  >} � 0   �}  �B  �|  �B  
 {*  u(  �#  "d  HN�,  mo P�.   ��  QM6  cmd R 6  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  gY6  8�W  hi6  P��  iy  h�� l�.  l�N  mR  |E�  pR  ��W  ry6  �~�  s�.  �*� t�.  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��.  �#�R  ��    #��  ��   #�  ��   #h  ��6  #I�  �y  @ �*  �z �(  �  	��  ��   	�\  �y  	�  ��,  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  ��,  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	�-  x E�   y F�   �{ Hp-  (T	�-  `e V�   x W�  y X�  z Y�    	�  [�-  �a	�.  = c�   F�  d�  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  o�.  ��  r
�.   iK  u�-  0��  x
�   XS�  {�.  `��  ~R   h��  ��   pu| ��/  x �,  �   �.  =    �}  X��/  v1 �E0   v2 �E0  dx ��  dy ��  �  �B  �k �B  tag �B  �W  ��  �o �K0  $��  �90  4SX  � 0  8d�  � 0  @��  �
�   H��  �R   P �/  �.  �z ��-  �	 0  2�  ��   ]  ��  �h  �B  �N  �B  
�K  �B  >} � 0   �/  �}  ��/  
K   �90  ��   �  o�  ��   ��  �0  �-  �  [0  =    �u  ��.  �z �{*  8�	�0  v1 �E0   v2 �E0  82  ��  Mp �$  [�  ��0   �  ��0   SX  � 0  (d�  � 0  0 0  [0  A{ �s0  4	T1  $x �   $y 	�  $dx 
�  $dy �  �o T1  )�  �  0 �  j1  =   =    (} �0  �  *�  %v  @292  @�  492   $x1 5�   $x2 6�   .]  8�  5]  9�  �� :�  ��  =�   �  @�   ��  C�  $�n  G?2  (9x  H?2  0�^  I?2  8 �0  B  >�  K�1  %�h  PR.3  s�  U.3   �H  V.3  $x1 X�   $x2 Y�   $gx \�  $gy ]�  $gz `�   $gzt a�  $�x  d�  (� f�  ,~�  i�  0t  k�  4.� l�   8�  p43  @	�  r�   H R2  w1  �h  tR2  �	|3  �c  �y   �O  �|3  �x  �
�3   B  �3  =    �  �3  =    I�  �G3  �	�3  �  ��    �  ��3   �3  �  ��3  &��	�4    ��   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  $top �	�4  '��  �	�  U'��  �	�  V'� �	�4  W'�  �	�  � �  �4  =   ? ��  ��3  	5  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�4  5  5  =    	S�  '5  
K   7L5  {�   U�  ~�   >	�5  �� @�*   s A
�   sx B�  sy C�   Nz EL5   	 6  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�5  
K   1M6  ��   ��  ��   �y  9,6  �   i6  =    y  y6  =    y  �6  =    �5  �6  =    hy ��*  (�		7  in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�.  �a  �
�   $ ��  ��6  ��	�7  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��7  ( 	7  �7  =    ޴  �7  	.L  &�7  �  	׮  )�7  	�  +�7  	�  ,�7  	�Q  .43  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7H8  �   	��  8H8  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�8  �3  	��  H�   	��  IE0  	��  K�   	a� L92  	w�  N�   	P{ O 0  	��  Q�   	��  R�8  g0  	��  T�   	�� U9  j1  	�}  W�   	u| X�0  	M�  Z�   	P�  [�0  	��  a�  	��  b�  	�  c�  	�p  e$  	�T  f�9  �6  	�a  j$  �   �9  =   � 	ը  l�9  $  �9  =   @ 	�p  m�9  	 �  p�  	p|  q$  	$Y  v�   	�K  y�   	g  {:  �4  	d�  |:  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   43  �:  =   =   / 	��  E�:  43  �:  =   / 	Ԁ  F�:  43  
;  =   =    	7� G�:  	�R  I�   	��  J43  	��  U�   (	P�  \G;  :;  	��  ]G;  	L�  ^G;  	ߵ  _G;  	�  aG;  	@�  92  	[�  �0  	 �  �0  	SX   0  	d�   0  	��  �   	_�   �   	��  "y  	��  %y  	'�  &y  	�]  (y  E2  <  =   � 	�P  *<  	ӯ  +)<  E2  	|  -;<  43  	��  .;<  	��  /;<  _<  o<  �   �    	��  ?2  �   Y<  	qY  "{<  	�  #{<  B  �<  =   ? 	��  %�<  	��  &�<  �  �<  =   � 	@Y  (�<  �  �<  =   ? 	V�  )�<  :3  =  =    	�h  =  	�  )=  :3  	�  :3  	�f  !�<  	r�  "�<  	��  %?2  	��  &?2  	׆  '�  	��  (�  	�  *�  	��  +�  	�  43  	��  �   	�_  �   	�_  �   	b  �  	t  �  	j�  "�,  	�  :�   	��  ;�   	��  <�   	�W  >43  	hn  @�  	U~  A�  	�  B�  	 �  C�  	%�  F�,  	�u  H�,  	z  I�,  	ʓ  C�  "  �>  =    	��  b>  �   �>  =    	��  c�>  	0K  d�   	?�  e�   �	?  x ��   y ��  dx ��  dy ��   ��  ��>  �5?  �p �
�.  ��  �
�0   �	d?  {q ��   ��  �y  d �	?   t�  �5?  d?  �?  =   � 	r �p?  	�T  ��?  d?  	l�  ��  	�  ��  	?k  ��  	�d  ��  	2~ �?  	��  �y  	��  ��  	k�  ��  	Z�  ��0  �0  @  =    	�v  �
@  	�v  ��   	"�  ��.  �  �,  �U  ?2  ��  ?2  t�  �   �  	�   .Y  
�  7Y  �  �h  �@  �.  *� �.  <i  �.  	G  y  	��  �   
K   ��@  )top  �G  �  �]  ��@   �	VA  ��  ��0   ��  ��@  O{  �
�   ��  �
�   iK  �VA   �-  ��  �A  \A  xA  =    	��  �hA  !K   �A  )up  �  �F  �S   FT  
�A  !K   �A  ��   �x  H�  ��  �H   ��  �A  H	�B  `e �   >}  0  L� �   $low �  $+�  �  (�Z !
�   ,r� "
�   0�f  #�A  4�f  $�A  8��  %y  <$tag &
�   @*� '�A  D �w )�A  �B  �B  =    �B  �  2�B  !K   �
C  ��   �s  z�  ��  �T  ܭ   gY  ��B  H�	�C  `e ��   *� �
C  >} � 0   �W  ��  (�}  ��  ,L� ��  0��  �y  4��  �
�   8$tag �
�   <��  �
�   @  w �C  �C  �C  =    �C  j�  �C   6  	��  My  	(h  N�   	l�  N�   	�  .y  	�  /y  	�  0y  	�  2y  	w�  8�  	�  9�  	�  :J  	�_  ;�   	��  >y  	�  Jy  	"�  R�  	t�  S�   	�w  T�   	؜  Y�   	q�  [y  	Ƚ  ^�  	�  _�   	�y  `�   	b�  c�   	+�  fy  	��  iy  	֘ l�   	�J  x�   	��  y�   	ks  �   	�  ��   	J�  ��   	�i  ��   	��  �y  	��  �y  	��  �y  	<� �y  	��  �y  	��  �y  	5�  �y  	<m  ��   	 K  ��   	�R  ��   	op  ��   	�m  ��   	D  ��   	X�  ��   	If  ��   	� ��   	��  �y  	�U  �y  	`  �y  	J�  �y  	��  �y  	� ��  �6  pF  =    	�  �`F  y  �F  =    	� �|F  "  �F  =   	 	,�  ��F  	R�  ��F  "  "  �F  =    	�u  ��F  	��  ��7  	�e  ��   �   G  =   � 	(�  ��F  	�  �y  ��  �  �v  �   n�  �   4�  �   *b �   ��  �C  *F  	Pif     *s>  (	`if     +�, {�vA     x       ��G  ,i }
�   r� n� -�vA     �H  - wA     �G  -wA     I  -
wA     I   +�� ^VvA     E       �UH  .Ye `UH  �� �� /�vA      I  DH  0Us  1�vA     0Us   �  +�� UUvA            ��H  2`e U$UH  U +c ILvA     	       ��H  2`e I"UH  U +3b :.vA            ��H  2`e :UH  U 3Yw .vA            �4�� �� V4�~ �~ -	4�s �s h4� � 7	 |L   &�  S#  D� �*  wA     ~      I ��  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �  
K   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
K   /  ��   [r  �4 #�  �   �X  5�  
K   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K&  
�   P�  =_  ��   R�  N�  ��  ��   �p  W�  
K   3�  ��   ({  ��  ğ   F]  8�  
K   Y@  ��   �c  |  ��  l  ��  �   
K   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {@  
K   ��  &�   �  º  GY  �f  ��   v�  ��  
K   �  GQ   ϼ  �  �_  X  &�  �b   
K   	Kf  � � ^�  �� e  2 8� ��  �  _�  �   t�  
 �   f  r  �  =   �' w  	��  1�  	]  4�  r  r  �  =   � �  	Zy  8�  �  �  =   =   � �  	��  ;�  Ʃ  QK   �       =       	�  W  �p  #3  9  @   S�  $L  R  ]  R    T}  %i  o    R   R    '	�  acv )'  ��  *@  ��  +]   �y -  �Y  6�  ��  :�  s�  <�   �H  =�  xz  >�   �  x @�  B    =    4  ,  =    
�	s  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x �,  
K   �	  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �  
K   �c#  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�	  (x	�#  �u z�	   � {	�   s |	�   � ~�  N�  c#  ��  �	�   ��  �	�     J]  �p#  �#  �#  =   � �^  ��#  �   $    �  �$  !K   �l'  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o   $  \	�(  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /y'  �(  �(  =   � ��  1�(  
K   p�)  �! 9& +! v( %# 0  B& @�! ��"  w#  	$  �-  S%  �)   0  @&  ��"    !0    m0    b-    �.    �$     /   @ %   � <"    U-    5'    	!  �]  ���+  `e �    x �f  y �f  z �f   ��  ��+  (cN  ��+  0Mp ��  8�u ��	  <� ��   @�H  ��+  Hr�  ��+  P��  ��+  X��  �f  `m�  �f  d��  �f  h  �f  l3F  �f  p8F  �f  t=F  �f  x��  ��   |*� �l'  �y� ��+  �s ��   ��� ��+  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  �+  ���  �   ���  	�   ��R  �-  �f�  �   �I}  s  ���  �+  � �)  Gx  ��+  >} �11   �}  �B  �|  �B  
 �+  �(  �#  "d  HN�-  mo P�/   ��  Q~7  cmd RQ7  �  Wf  (_  Yf   #_  [f  $bob ]f  (�  a�   ,�[  b�   0sb  d�   4d]  g�7  8�W  h�7  P��  iy  h�� l�/  l�N  m�  |E�  p�  ��W  r�7  �~�  s�/  �*� t�/  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��/  �#�R  ��    #��  ��   #�  ��   #h  ��7  #I�  �y  @ �+  �z �)  �  	��  ��   	�\  �y  	�  �
.  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  ��-  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	�.  x Ef   y Ff   �{ H�.  (T	/  `e V    x Wf  y Xf  z Yf    	�  [�.  �a	�/  = cf   F�  df  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  o�/  ��  r
�/   iK  u/  0��  x
�   XS�  {�/  `��  ~R   h��  ��   pu| ��0  x �-  �   0  =    �}  X��0  v1 �v1   v2 �v1  dx �f  dy �f  �  �B  �k �B  tag �B  �W  �  �o �|1  $��  �j1  4SX  �11  8d�  �11  @��  �
�   H��  �R   P �0  0  �z �/  �	11  2�  �f   ]  �f  �h  �B  �N  �B  
�K  �B  >} �11   �0  �}  ��0  
K   �j1  ��   �  o�  ��   ��  �C1  �.  f  �1  =    �u  �0  �z ��+  8�	2  v1 �v1   v2 �v1  82  �f  Mp ��  [�  �2   �  �2   SX  �11  (d�  �11  0 71  �1  A{ ��1  4	�2  $x f   $y 	f  $dx 
f  $dy f  �o �2  )�    0 f  �2  =   =    (} ,2  �  *�  %v  @2j3  @�  4j3   $x1 5�   $x2 6�   .]  8f  5]  9f  �� :f  ��  =�   �  @f   ��  Cf  $�n  Gp3  (9x  Hp3  0�^  Ip3  8  2  B  >�  K�2  %�h  PR_4  s�  U_4   �H  V_4  $x1 X�   $x2 Y�   $gx \f  $gy ]f  $gz `f   $gzt af  $�x  df  (� ff  ,~�  if  0t  kf  4.� l�   8�  pe4  @	�  r�   H �3  �2  �h  t�3  �	�4  �c  �y   �O  ��4  �x  �
�4   B  �4  =    �  �4  =    I�  �x4  �	5  �  ��    �  �5   �4  �  ��4  &��	�5    �f   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  $top �	�5  '��  �	�  U'��  �	�  V'� �	�5  W'�  �	�  � �  �5  =   ? ��  �5  	46  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�5  46  P6  =    	S�  '@6  
K   7}6  {�   U�  ~�   >	�6  �� @�+   s A
�   sx Bf  sy Cf   Nz E}6   	Q7  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�6  
K   1~7  ��   ��  ��   �y  9]7  
K   @�7  el �l �l  �   �7  =    y  �7  =    y  �7  =    �6  �7  =    hy ��+  (�	[8  in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�/  �a  �
�   $ ��  ��7  ��	 9  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  � 9  ( [8  9  =    ޴  �g8  	.L  &(9  f  	׮  )(9  	�  +(9  	�  ,(9  	�Q  .e4  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�9  �   	��  8�9  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�9  5  	��  H�   	��  Iv1  	��  K�   	a� Lj3  	w�  N�   	P{ O11  	��  Q�   	��  RN:  �1  	��  T�   	�� Ul:  �2  	�}  W�   	u| X2  	M�  Z�   	P�  [2  	��  af  	��  bf  	�  cf  	�p  e�  	�T  f�:  �7  	�a  j�  �   ;  =   � 	ը  l�:  �  ;  =   @ 	�p  m;  	 �  pf  	p|  q�  	$Y  v�   	�K  y�   	g  {f;  �5  	d�  |f;  	��   f  		�  !f  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +f  	`�  ,f  	A�  -f  	��  /�   	��  1�   	P�  2�   e4  <  =   =   / 	��  E<  e4  :<  =   / 	Ԁ  F*<  e4  \<  =   =    	7� GF<  	�R  I�   	��  Je4  	��  U�   (	P�  \�<  �<  	��  ]�<  	L�  ^�<  	ߵ  _�<  	�  a�<  	@�  j3  	[�  2  	 �  2  	SX  11  	d�  11  	��  �   	_�   �   	��  "y  	��  %y  	'�  &y  	�]  (y  v3  c=  =   � 	�P  *S=  	ӯ  +{=  v3  	|  -�=  e4  	��  .�=  	��  /�=  �=  �=  �   �    	��  p3  �   �=  	qY  "�=  	�  #�=  B  >  =   ? 	��  %�=  	��  &�=  f  *>  =   � 	@Y  (>  f  G>  =   ? 	V�  )6>  k4  c>  =    	�h  S>  	�  {>  k4  	�  k4  	�f  !�=  	r�  "�=  	��  %p3  	��  &p3  	׆  'f  	��  (f  	�  *f  	��  +f  	�  e4  	��  �   	�_  �   	�_  �   	b  f  	t  f  	j�  "�-  	�  :�   	��  ;�   	��  <�   	�W  >e4  	hn  @f  	U~  Af  	�  Bf  	 �  Cf  	%�  F�-  	�u  H�-  	z  I�-  	ʓ  C   s  �?  =    	��  b�?  �   �?  =    	��  c�?  	0K  d�   	?�  e�   �	Y@  x �f   y �f  dx �f  dy �f   ��  �!@  ��@  �p �
�/  ��  �
2   �	�@  {q �f   ��  �y  d �	e@   t�  ��@  �@  �@  =   � 	r ��@  	�T  ��@  �@  	l�  �f  	�  �f  	?k  �f  	�d  �f  	2~ �Y@  	��  �y  	��  �f  	k�  �f  	Z�  �2  2  lA  =    	�v  �\A  	�v  ��   	"�  ��/  �  �-  �U  p3  ��  p3  t�  �   �  	�   .Y  
f  7Y  f  �h  �A  �/  *� �/  <i  �/  	G  y  	��  �   
K   �QB  )top  �G  �  �]  �0B   �	�B  ��  �2   ��  �QB  O{  �
�   ��  �
�   iK  ��B   /  ��  �]B  �B  �B  =    	��  ��B  !K   �B  )up  �  �F  �S   FT  
�B  !K   8C  ��   �x  H�  ��  �H   ��  
C  H	�C  `e     >} 11  L� f   $low f  $+�  f  (�Z !
�   ,r� "
�   0�f  #�B  4�f  $�B  8��  %y  <$tag &
�   @*� '8C  D �w )EC  D  D  =    �C  �  2D  !K   �\D  ��   �s  z�  ��  �T  ܭ   gY  �(D  H�	 E  `e �    *� �\D  >} �11   �W  �f  (�}  �f  ,L� �f  0��  �y  4��  �
�   8$tag �
�   <��  �
�   @  w �iD  E  E  =     E  j�  E  Q7  	��  My  	(h  N�   	l�  N�   	�  .y  	�  /y  	�  0y  	�  2y  	w�  8  	�  9�  	�  :�  	�_  ;�   	��  >y  	�  Jy  	"�  R�  	t�  S�   	�w  T�   	؜  Y�   	q�  [y  	Ƚ  ^�  	�  _�   	�y  `�   	b�  c�   	+�  fy  	��  iy  	֘ l�   	�J  x�   	��  y�   	ks  �   	�  ��   	J�  ��   	�i  ��   	��  �y  	��  �y  	��  �y  	<� �y  	��  �y  	��  �y  	5�  �y  	<m  ��   	 K  ��   	�R  ��   	op  ��   	�m  ��   	D  ��   	X�  ��   	If  ��   	� ��   	��  �y  	�U  �y  	`  �y  	J�  �y  	��  �y  	� ��  �7  �G  =    	�  ��G  y  �G  =    	� ��G  s  �G  =   	 	,�  ��G  	R�  �H  s  s  (H  =    	�u  �H  	��  �9  	�e  ��   �   ]H  =   � 	(�  �LH  	�  �y  ��  �  �v  �   n�  �   4�  �   *b �   ��  0E  *�� ,
y  	xif     +�� ��yA     �      ��I  ,�R  ��:  م υ -cmd �0E  X� N� .� ��  ݆ ׆ /�yA     �I  LI  0U�U 1�yA     NJ  2zA     �J  qI  0Us  2zA     7L  �I  0Us  2�zA     CL  �I  0Us  3�zA     OL  0Us   +� ��xA     �       �NJ  ,�R  ��:  0� *� .Mp ��  ~� |� .� ��  �� �� 2�xA     OL  (J  0Us  2)yA     �J  @J  0Us  1NyA     [L   +΀ �TxA     �       ��J  ,�R  ��:  Ї Ƈ -cmd �0E  O� E� 2�xA     K  �J  0Us  2�xA     K  �J  0Us  4�xA     gL  0T�  5� FK  6�R  F�:  7Mp H
�   8bob If   +(� 4wA     B       ��K  ,�R  5�:  Ԉ Έ ,Mp 6�  (�  � ,��  7f  �� �� 23wA     sL  }K  0U|  3IwA     sL  0U|   9�J  UwA     �       �7L  :�J  � ۉ ;�J  ;�J  <�J  �wA     �       L  :�J  /� -� =�wA     �       ;�J  >�J  T� R� 1�wA     sL    1hwA     sL  1wwA     sL   ?Q Q A	?�o �o �?�u �u O?Ef Ef x?�e �e s	?d  d  
"	 �G   ��  S#  v� �*  �{A           � �  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �  
K   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
K   /  ��   [r  �4 #�  �   �X  5�  
K   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K&  
�   P�  =_  ��   R�  N�  ��  ��   �p  W�  
K   3�  ��   ({  ��  ğ   F]  8�  
K   Y@  ��   �c  |  ��  l  ��  �   
K   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {@  
K   ��  &�   �  º  GY  �f  ��   v�  ��  
K   �  GQ   ϼ  �  �_  X  &�  �b   t�  	 �     
K   
M  �L  M M �L   	�  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4M  �  	D  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�  D  `  =    	S�  'P  !  }  =   �' l  	��  1}  	]  4�  !  !  �  =   � �  	Zy  8�  �  �  =   =   � �  	��  ;�  Ʃ  QK   �  �    =     �  	�  W  �p  #(  .  5   S�  $A  G  R  R    T}  %^  d  t  R   R    '	�  acv )  ��  *5  ��  +R   �y -t  �Y  6�  ��  :�  s�  <�   �H  =�  xz  >�   �  x @�  
K   R
  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �  
K   ��#  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u^
  (x	_$  �u zR
   � {	�   s |	�   � ~�  N�  �#  ��  �	�   ��  �	�     J]  ��#  _$  }$  =   � �^  �l$  �   �$    �  ��$  !K   ��'  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �$  \	H)  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /�'  H)  e)  =   � ��  1U)  
K   7�)  {�   U�  ~�   >	�)  �� @�)   s A
�   "sx B  "sy C   _$  Nz E�)  B  �)  =    4  *  =    
�	H*  "x �B   "y �B  Mp �B  *� �B  ޽  �B   ~x �*  �]  ��*,  `e ��   "x �  "y �  "z �   ��  �*,  (cN  �*,  0Mp ��  8�u �R
  <� ��   @�H  �*,  Hr�  �*,  P��  �e,  X��  �  `m�  �  d��  �  h  �  l3F  �  p8F  �  t=F  �  x��  ��   |*� ��'  �y� �k,  �s ��   ��� ��)  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  *,  ���  �   ���  	�   ��R  K.  �f�  �   �I}  H*  ���  *,  � T*  Gx  �e,  >} �M3   �}  �B  �|  �B  
 0,  H)  #d  HNK.  "mo P�.   ��  Q�.  "cmd R�  �  W  (_  Y   #_  [  $"bob ]  (�  a�   ,�[  b�   0sb  d�   4d]  g�.  8�W  h�.  P��  iy  h�� l�.  l�N  m�  |E�  p�  ��W  r�.  �~�  s�.  �*� t�.  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��.  �$�R  ��    $��  ��   $�  ��   $h  ��.  $I�  �y  @ q,  �z T*  �  
K   1�.  ��   ��  ��   �y  9d.  Q.  �   �.  =    y  �.  =    �   �.  =    y  �.  =    �)  �.  =    hy �q,  (�	W/  "in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�.  �a  �
�   $ ��  ��.  ��	�/  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��/  ( W/  0  =    ޴  �c/  	��  ��   	�\  �y  	�  �<0  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  �^.  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	�0  "x E   "y F   �{ H�0  (T	71  `e V�   "x W  "y X  "z Y    	�  [�0  �a	2  = c   F�  d  �~ eB  h�  fB  
t�  gB  �k hB  "tag iB  �N  l
�   ��  o�.  ��  r
�.   iK  u71  0��  x
�   XS�  {�.  `��  ~R   h��  ��   pu| ��2  x �}  X��2  "v1 ��3   "v2 ��3  "dx �  "dy �  �  �B  �k �B  "tag �B  �W  ��)  �o ��3  $��  ��3  4SX  �M3  8d�  �M3  @��  �
�   H��  �R   P �2  2  �z �C1  �	M3  2�  �   ]  �  �h  �B  �N  �B  
�K  �B  >} �M3   �2  �}  ��2  
K   ��3  ��   �  o�  ��   ��  �_3  �0    �3  =    �u  �2  �z �0,  8�	04  "v1 ��3   "v2 ��3  82  �  Mp ��  [�  �04   �  �64   SX  �M3  (d�  �M3  0 S3  �3  A{ ��3  4	�4  %x    %y 	  %dx 
  %dy   �o �4  )�  �)  0   �4  =   =    (} H4  �  *�  &v  @2�5  @�  4�5   %x1 5�   %x2 6�   .]  8  5]  9  �� :  ��  =�   �  @   ��  C  $�n  G�5  (9x  H�5  0�^  I�5  8 <4  B  >�  K�4  &�h  PR{6  s�  U{6   �H  V{6  %x1 X�   %x2 Y�   %gx \  %gy ]  %gz `   %gzt a  $�x  d  (� f  ,~�  i  0t  k  4.� l�   8�  p�6  @	�  r�   H �5  �4  �h  t�5  �	�6  �c  �y   �O  ��6  �x  �
�6   B  �6  =    �  �6  =    I�  ��6  �	7  �  ��    �  �7   �6  �  ��6  '��	�7    �   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  %top �	�7  (��  �	�  U(��  �	�  V(� �	�7  W(�  �	�  � �  �7  =   ? ��  �07  	.L  &8    	׮  )8  	�  +8  	�  ,8  	�Q  .�6  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7v8  �   	��  8v8  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�8  #7  	��  H�   	��  I�3  	��  K�   	a� L�5  	w�  N�   	P{ OM3  	��  Q�   	��  R*9  �3  	��  T�   	�� UH9  �4  	�}  W�   	u| X64  	M�  Z�   	P�  [04  	��  a  	��  b  	�  c  	�p  e�  	�T  f�9  �.  	�a  j�  �   �9  =   � 	ը  l�9  �  �9  =   @ 	�p  m�9  	 �  p  	p|  q�  	$Y  v�   	�K  y�   	g  {B:  �7  	d�  |B:  	��     		�  !  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +  	`�  ,  	A�  -  	��  /�   	��  1�   	P�  2�   �6  �:  =   =   / 	��  E�:  �6  ;  =   / 	Ԁ  F;  �6  8;  =   =    	7� G";  	�R  I�   	��  J�6  	��  U�   	P�  \�  	��  ]�  	L�  ^�  	ߵ  _�  	�  a�  	��  �5  �   �;  �;  �;  �   �    	qY  "�;  	�  #�;  B  �;  =   ? 	��  %�;  	��  &�;    #<  =   � 	@Y  (<    @<  =   ? 	V�  )/<  �6  \<  =    	�h  L<  	�  t<  �6  	�  �6  	�f  !�;  	r�  "�;  	��  %�5  	��  &�5  	׆  '  	��  (  	�  *  	��  +  �  	��  My  	(h  N�   	l�  N�   	�  .y  	�  /y  	�  0y  	�  2y  	w�  8  	�  9�  	�  :�  	�_  ;�   	��  >y  	�  Jy  	"�  R�  	t�  S�   	�w  T�   	؜  Y�   	q�  [y  	Ƚ  ^�  	�  _�   	�y  `�   	b�  c�   	+�  fy  	��  iy  	֘ l�   	�J  x�   	��  y�   	ks  �   	�  ��   	J�  ��   	�i  ��   	��  �y  	��  �y  	��  �y  	<� �y  	��  �y  	��  �y  	5�  �y  	<m  ��   	 K  ��   	�R  ��   	op  ��   	�m  ��   	D  ��   	X�  ��   	If  ��   	� ��   	��  �y  	�U  �y  	`  �y  	J�  �y  	��  �y  	� ��  �.  x?  =    	�  �h?  y  �?  =    	� ��?  H*  �?  =   	 	,�  ��?  	R�  ��?  H*  H*  �?  =    	�u  ��?  	��  �0  	�e  ��   �   @  =   � 	(�  �@  	�  �y  ��  �  �v  �   n�  �   4�  �   *b �   ��  �<  )@�  (	�5  	Ъf     )[�  )
04  	�if     ) �  *
64  	�jf     )SX  +M3  	�if     )d�  ,M3  	Ȫf     �5  �@  =   � )�P  .�@  	�jf     )ӯ  /#A  	��f     �5  I	MA  �~ K	�    r�  L	�    1� N)A  )ف ToA  	�if     MA  MA  �A  =    )\� UuA  	�if     �   �A  =   =    *D� f�A  	�ae     +f� !�A     �       �rB  ,~ !�   �� w� -bsp #H9  � � .<p $
�   P� H� /(�A     rB  0U�A     cG  KB  1Qs  2i�A     �A  3y�A     FC  1Uv4$s "  +�� �>A     �       �FC  4num ��   �� �� .r� ��   � � .��  ��5  3� +� -sub �*9  �� �� 0\A     oG  
C  1U	��B     1Ts  2�A     {G  2�A     {G  2�A     �G  3�A     �D  1UsH  5%� v	y  ~A     "      ��D  ,�� v8  �� �� .~� x�   
� � 6�� y�   .=� z�   1� -� -x1 |  i� g� -y1 }  �� �� -x2 ~  � � -y2   � � .'Y  ��  A� ;� .p� ��  �� �� .Z� ��  �  � .Y� ��  M� ?� .' �oA  �� � -sx1 ��   1� /� -sx2 ��   X� T� 2�~A     �G  3�~A     �G  1Uv 1T|   7ρ �
}A           ��E  8��  ��5  �� �� 9x1 ��   >� :� 9x2 ��   |� t� .'Y   �  � ܑ .p� �  9� /� .Z� �  �� �� .Y� �  +� � :�� [~A     :�� W~A     2$}A     �G  24}A     �G  /~A     �E  /~A     sF   ;� ��|A     -       �7�� ��|A     Y       �sF  8�~ ��   �� �� 8r�  ��    � �� <' �oA  �� �� 0�|A     �G  PF  1U�U 2�|A     �G  =�|A     �G  1T�T  7�� a�{A     �       �IG  8�~ b	�   � �� 8r�  c	�   b� \� <�H  eoA  �� �� <' foA  J� @� >)o �Y|A     0�{A     �G  G  1Uv 1T|  0|A     �G  'G  1Uv  2<|A     �G  3U|A     �G  1T|   ;� =�{A            �?� � g?��  ��  7?M� M� ??O� O� 3?w� w� s?_� _� 3 <`   @�  S#  � �*  ��A     U      6( ��  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �  	"|  *y  	��  +y  	I�  ,y  	�a  -y   	R  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�  d  
K   	"�  ��  WH  �~  �O  �m  ��   �  ��  ��  	 
K   
�  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  
(�  
K   
/.  ��   [r  �4 #�  �   �X  
5  
K   
:�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  
K:  
�   
P�  =_  ��   R�  N�  ��  ��   �p  
W�  =� �  ��  .)  ^�  2�   }�  7�  �� ;K    	Z  r�  o   .� $�  O� )�   i  i  �    �  Z  �  i   u  1   �  i  K   R   1    �  ��  ,)  �  �  oS  '�  dS  ()*  � +
*   � ,i  @�  -
�   >z .
�   �  /R   �H  3:    �   :  =    �  	�� 7:  	�� 8K   
K   3  ��   ({  ��  ğ   F]  8X  
K   Y�  ��   �c  |  ��  l  ��  �   
K   k  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {�  
K   �T  &�   �  º  GY  �f  ��   v�  �!  
K   ��  GQ   ϼ  �  �_  X  &�  �b   t�   �   �  �  �  =   �' �  	��  1�  	]  4�  �  �  �  =   � �  	Zy  8�  �    =   =   �    	��  ;  Ʃ  QK   '  3  I  =     8  	�  WI  �p  #f  l  s   S�  $  �  �  R    T}  %�  �  �  R   R    '	�  acv )Z  ��  *s  ��  +�   �y -�  �Y  6�  ��  :-  s�  <-   �H  =-  xz  >�   �  x @�  B  O  =    4  _  =    
�	�  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x �_  
K     @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  
K   ��%  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u  (x	&   �u z    � {	�    s |	�    � ~�   N�  �%   ��  �	�    ��  �	�     J]  ��%  &  .&  =   � !�^  �&  �   F&  " !�  �;&  #K   ��)  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  S&  \	�*   �Y  	�     *O  	�    ��  	�    �  	�    b�  	�    ��  	�    �  	�    +�  	�    Zp  	�     o�   	�   $ m�  !	�   ( 4�  "	�   , �  #	�   0 �  $	�   4 ��  %	�   8 L� &	�   < ��  '	�   @   (	�   D ��  )	�   H \q *	�   L z�  +	�   P �  ,	�   T /�  -	�   X ʤ  /�)  �*  +  =   � !��  1+  �]  ���,  `e �3   x ��  y ��  z ��   ��  ��,  (cN  ��,  0Mp �'  8�u �  <� ��   @�H  ��,  Hr�  ��,  P��  �4-  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� ��)  �y� �:-  �s ��   ��� �@-  ��  ��   ��  ��   �ʺ  ��   ��l  ��   �  �  �,  � ��  �   � ��  	�   � �R   /  � f�  �   � I}  �  � ��  �,  � #+  Gx  �4-  >} �!3   �}  �B  �|  �B  
 �,  �*  &  $d  HN /  mo P�1   ��  Q�8  cmd RR  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g�8  8�W  h�8  P��  iy  h�� l�1  l�N  m  |E�  p  ��W  r9  �~�  s�1  �*� t�1  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��1  �%�R  ��    %��  ��   %�  ��   %h  �9  %I�  �y  @ F-  �z #+  	��  ��   	�\  �y  	�  �W/  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  ��  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   (	90  ��  B      B  Vd  !B  �  "B  �� #90   �   I0  =    � %�/  (	y0  � *�   �� +�   � ,U0  G /y0  C	�0  x E�   y F�   �{ H�0  (T	�0  `e V3   x W�  y X�  z Y�    	�  [�0  �a	�1  = c�   F�  d�  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  o�1  ��  r
�1   iK  u�0  0��  x
�   XS�  {�1  `��  ~R   h��  ��   pu| ��2  x &/  �   �1  =    �}  X��2  v1 �f3   v2 �f3  dx ��  dy ��  �  �B  �k �B  tag �B  �W  �?  �o �l3  $��  �Z3  4SX  �!3  8d�  �!3  @��  �
�   H��  �R   P �2  �1  �z �1  �	!3  2�  ��   ]  ��  �h  �B  �N  �B  
�K  �B  >} �!3   �2  �}  ��2  
K   �Z3  ��   �  o�  ��   ��  �33  �0  �  |3  =    �u  ��1  �z ��,  8�	4  v1 �f3   v2 �f3  82  ��  Mp �'  [�  �4   �  �
4   SX  �!3  (d�  �!3  0 '3  |3  A{ ��3  4	u4  &x �   &y 	�  &dx 
�  &dy �   �o u4   )�  O  0 �  �4  =   =    (} 4  �  *�  'v  @2Z5   @�  4Z5   &x1 5�   &x2 6�    .]  8�   5]  9�   �� :�   ��  =�    �  @�    ��  C�  $ �n  G`5  ( 9x  H`5  0 �^  I`5  8 4  B  >�  K�4  '�h  PRO6   s�  UO6    �H  VO6  &x1 X�   &x2 Y�   &gx \�  &gy ]�  &gz `�   &gzt a�  $ �x  d�  ( � f�  , ~�  i�  0 t  k�  4 .� l�   8 �  pU6  @ 	�  r�   H s5  �4  �h  ts5  �	�6   �c  �y    �O  ��6   �x  �
�6   B  �6  =    �  �6  =    I�  �h6  �	�6   �  ��     �  ��6   �6  �  ��6  (��	�7     ��    �  �	�    t�  �	�    ��  �	�    /�  �	�    �  �	�  &top �	�7  )��  �	�  U)��  �	�  V)� �	�7  W)�  �	�  � �  �7  =   ? ��  �7  	$8  ~�  T   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�7  $8  @8  =    	S�  '08  
K   7m8  {�   U�  ~�   >	�8  �� @@-   s A
�   sx B�  sy C�   Nz Em8  
K   1�8  ��   ��  ��   �y  9�8  �   �8  =    y  9  =    y  9  =    �8  "9  =    hy �F-  (�	�9  in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�1  �a  �
�   $ ��  �.9  ��	7:  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  �7:  ( �9  G:  =    ޴  ��9  	.L  &_:  �  	׮  )_:  	�  +_:  	�  ,_:  	�Q  .U6  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�:  �   	��  8�:  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F;  �6  	��  H�   	��  If3  	��  K�   	a� LZ5  	w�  N�   	P{ O!3  	��  Q�   	��  R�;  �3  	��  T�   	�� U�;  �4  	�}  W�   	u| X
4  	M�  Z�   	P�  [4  	��  a�  	��  b�  	�  c�  	�p  e'  	�T  f<  "9  	�a  j'  �   8<  =   � 	ը  l'<  '  U<  =   @ 	�p  mD<  	 �  p�  	p|  q'  	$Y  v�   	�K  y�   	g  {�<  �7  	d�  |�<  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   U6  U=  =   =   / 	��  E?=  U6  q=  =   / 	Ԁ  Fa=  U6  �=  =   =    	7� G}=  	�R  I�   	��  JU6  	��  U�   	P�  \^  	��  ]^  	L�  ^^  	ߵ  _^  	�  a^  	@�  Z5  	[�  4  	 �  
4  	SX  !3  	d�  !3  	��  �   	_�   �   	��  "y  	��  %y  	'�  &y  	�]  (y  f5  �>  =   � 	�P  *�>  	ӯ  +�>  f5  	|  -�>  U6  	��  .�>  	��  /�>  �>  �>  �   �    	��  `5  �   �>  	qY  "�>  	�  #�>  B  2?  =   ? 	��  %!?  	��  &!?  �  Z?  =   � 	@Y  (J?  �  w?  =   ? 	V�  )f?  [6  �?  =    	�h  �?  	�  �?  [6  	�  [6  	�f  !!?  	r�  "!?  	��  %`5  	��  &`5  	׆  '�  	��  (�  	�  *�  	��  +�  	�  U6  	��  �   	�_  �   	�_  �   	b  �  	t  �  	j�  "�  	�  :�   	��  ;�   	��  <�   	�W  >U6  	hn  @�  	U~  A�  	�  B�  	 �  C�  	%�  F�  	�u  H�  	z  I�  	ʓ   C3  �  A  =    	��   bA  �   -A  =    	��   cA  	0K   d�   	?�   e�    �	�A  x  ��   y  ��  dx  ��  dy  ��   ��   �QA   ��A  �p  �
�1  ��   �

4    �	�A  {q  ��   ��   �y  d  �	�A   t�   ��A  �A  B  =   � 	r  ��A  	�T   �B  �A  	l�   ��  	�   ��  	?k   ��  	�d   ��  	2~  ��A  	��   �y  	��   ��  	k�   ��  	Z�   �
4  
4  �B  =    	�v   ��B  	�v   ��   	"�   ��1  !�   �  !�U   `5  !��   `5  !t�   �   !�   	�   !.Y   
�  !7Y   �  !�h   (C  �1  !*�  �1  !<i   �1  	G  !y  	��  !�   �   pC  =    
K   !��C  *top  �G  �  �]  !�pC   !�	�C  ��  !�
4   ��  !��C  O{  !�
�   ��  !�
�   iK  !��C   �0  ��  !��C  �C  
D  =    	��  !��C  #K   !=D  *up  �  �F  �S   FT  !
D  #K   !xD  ��   �x  H�  ��  �H   ��  !JD  H!	8E   `e !3    >} !!3   L� !�   &low !�  $ +� ! �  ( �Z !!
�   , r� !"
�   0 �f  !#=D  4 �f  !$=D  8 ��  !%y  <&tag !&
�   @ *� !'xD  D �w !)�D  UE  UE  =    8E  !�  !2EE  #K   !��E  ��   �s  z�  ��  �T  ܭ   gY  !�hE  H!�	@F   `e !�3    *� !��E   >} !�!3    �W  !��  ( �}  !��  , L� !��  0 ��  !�y  4 ��  !�
�   8&tag !�
�   < ��  !�
�   @  w !��E  ]F  ]F  =    @F  !j�  !MF  R  	��  "My  	(h  "N�   	l�  "N�   	�  #.y  	�  #/y  	�  #0y  	�  #2y  	w�  #8.  	�  #9�  	�  #:�  	�_  #;�   	��  #>y  	�  #Jy  	"�  #R�  	t�  #S�   	�w  #T�   	؜  #Y�   	q�  #[y  	Ƚ  #^�  	�  #_�   	�y  #`�   	b�  #c�   	+�  #fy  	��  #iy  	֘ #l�   	�J  #x�   	��  #y�   	ks  #�   	�  #��   	J�  #��   	�i  #��   	��  #�y  	��  #�y  	��  #�y  	<� #�y  	��  #�y  	��  #�y  	5�  #�y  	<m  #��   	 K  #��   	�R  #��   	op  #��   	�m  #��   	D  #��   	X�  #��   	If  #��   	� #��   	��  #�y  	�U  #�y  	`  #�y  	J�  #�y  	��  #�y  	� #�  "9  I  =    	�  #��H  y  I  =    	� #�I  �  :I  =   	 	,�  #�*I  	R�  #�RI  �  �  hI  =    	�u  #�XI  	��  #�G:  	�e  #��   �   �I  =   � 	(�  #��I  	�  #�y  !��  #  !�v  #�   !n�  #�   !4�  #�   !*b #�   !��  #pF  	- $�   	_  $ �   
;	fJ  C� =B   � >B  .� ?B  �� @B  �  AB   � BJ   J	�J  � L*   "� M�   ��  NB    OB  �� P�   Â QB  ;� R�J   fJ  �J  =     O� SrJ  Y	$K  C� ^B   � _B  .� `
�    ك a�J  R� h<K  ۄ (j�K  � m
*   ��  nB    oB  
�8 s�   �H  w�K  Â {B  ;� |�K   0K  $K  �K  =     +�:  �	��f     ,E� ��   	P�f     ,� ��   	 �f     ,�� ��   	(�f     ,#� ��   	h�f     ,8� ��   	��f     +�:  �	��f     +�:  �	$�f     +�:  �	تf     ,�� ��   	�f     ,�� ��L  	8�f     �K  ,�� ��L  	H�f     ,4� ��:  	`�f     +S:  �	0�f     ,�� ��:  	�f     ,� �M  	@�f     `5  ,{� �)M  	�f     /M  4  ,� �
KM  	�f     �  +�:  �	��f     +�:  �	x�f     +e:  �
	X�f     +q:  �
	�f     +}:  �
	 �f     +�:  �	p�f     -K� �   	�f     -�� �   	�f     -N� �   	��f     .�{  x�A     }      ��O  /C� "�   ̖ Ȗ /� #�   � � /� $�   B� <� 0i &�   �� �� 0j '�   :� 4� 1k (�   /�O  )�   �� �� /P{  +�K  � � 0th ,�O  � � 0sf -�6  5� 3� 2��A     �_  �N  3T13Q0 2.�A     �_  O  3T8 2;�A     �_  .O  3Us  2M�A     �_  JO  3T13Q0 2�A     �_  aO  3T8 2�A     �_  yO  3Us  2+�A     �_  �O  3T13Q0 2֍A     �_  �O  3T8 4�A     �_   3  5w! �   R�A     &       �EP  6�  �   ^� X� 0i 	
�   �� �� 2]�A     EP  #P  3Uv  7r�A     �_  3U	��B     3Tv   8e~ ��   P  9� �%�   :P{  ��K  1key �	�    5) ��   ��A     B       �Q  6� ��   �� �� 0i �
�   M� K� ;�� �
`C  �W2ʊA     �_  �P  3Uv  7�A     �_  3U	��B     3T�W  .ƃ ���A     1       ��Q  <��A     �S  2��A     �_  XQ  3U. <��A     %S  2��A     �_  }Q  3U. <��A     R  2��A     �_  �Q  3U. 4��A     �Q   .�� �k�A             �R  /�O  �	�   r� p� 2v�A     �_  R  3U	��B      7��A     �_  3T1  .΂ �w�A     �       �S  0i �
�   �� �� /.� �S  � � 2��A     �_  }R  3U	�WB      2��A     �_  �R  3U	I�B      2��A     �_  �R  3T13Qs  2މA     �_  �R  3T13Qs  2��A     �_  �R  3T13Qs  2�A     �_  S  3U. 70�A     �_  3T8  I0  .l� y�A     b       ��S  0i {
�   ?� 7� 2 �A     �_  vS  3U	��B      22�A     �_  �S  3U	�XB      7\�A     �_  3T13Q0  .�� ���A           �[Z  /�N  �[Z  �� �� /P{  ��K  � � /�� �aZ   � � /.� �gZ  I� C� 0i ��   �� �� 0j ��   �� u� /Ԅ ��:  m� e� /f� ��:  Ϡ ɠ /� ��:  � � ;� �`C  ��/� ��   V� R� /̈́ ��   �� �� /�� ��:  Ρ ʡ / ��   � � /� ��   .� ,� /82  ��   U� Q� /�� ��   �� �� /�� ��   � ޢ /)� ��   � � /6� ��   C� ?� /\� ��:  �� y� /�� ��   �� �� /�� ��   M� G� /�� ��   �� �� =mZ  r�A      r�A     �       qHV  >r�A     �       ?{Z  � � ?�Z  D� @� ?�Z  ~� z� 2��A     �_  9V  3T13Qv  <A     �_    2�A     �_  lV  3U	0�B     3T1 2:�A     �_  �V  3U| 2$3T13Qv  2Z�A     �_  �V  3U��3Tsx3Q9 2d�A     �_  �V  3U�� 2{�A     �_  �V  3U	0�B      2��A     �_  W  3U	7�B     3T1 2��A     �_  0W  3U	7�B      <��A     `  2��A     �_  \W  3U	@�B      2τA     �_  �W  3U	@�B     3T1 2ބA     �_  �W  3U	@�B      <�A     `  2�A     �_  �W  3Us 3$3T13Q0 24�A     �_  �W  3T13Q0 2T�A     �_  X  3T13Q0 2t�A     �_  $X  3T13Q0 2��A     �_  @X  3T13Q0 2��A     �_  \X  3T13Q0 2ԅA     �_  xX  3T13Q0 2�A     �_  �X  3U	�WB      2�A     �_  �X  3U	I�B      < �A     `  22�A     �_  �X  3U[ 2H�A     �_  �X  3U  2Z�A     �_  Y  3U] 2l�A     �_  "Y  3U8 2��A     �_  :Y  3U. 2�A     �_  YY  3U	O�B      2#�A     �_  uY  3T13Q0 2��A     �_  �Y  3U	u�B     3T}  2чA     �_  �Y  3T13Q0 2�A     �_  �Y  3T13Q0 2�A     �_  �Y  3U�� 2�A     �_  Z  3U	7�B      2-�A     �_  *Z  3U	@�B      2B�A     =[  BZ  3Us 7W�A     �_  3T13Q0  �J  fJ  $K  @b� ��Z  :�� ��L  1i �	�   1key �	�    5�� �  ��A     n       �=[  Atex ��   ̥ ¥ Acol ��   B� >� /�O  �
�   �� �� 0ofs �
�   �� �� 2΃A     �_  /[  3T8 <�A     �\   .[� &�A     �      ��\  6�� &�   �� �� /P{  (�K  � � ;Â )�  ��/.� *gZ  A� 7� /x� +S  ب ֨ 0x ,�   	� �� 0x1 -�   �� �� 0x2 .�   ͩ ǩ 0i /�   )� #� /у 0`5  v� t� /-� 1/M  �� �� 2r�A     �_  W\  3T13Q�� 2��A     �_  n\  3T8 2&�A     `  �\  3U	��B     3Ts  2a�A     �_  �\  3U	�B     3T~  <{�A     �_   B$� ��A           �4^  C�� ��   Ī �� D�� ��  � � DP{  ��K  a� _� D.� �gZ  �� �� Dx� �S  %� #� Ex ��   P� H� Ex1 ��   ¬ �� Ex2 ��   � � Ei ��   '� � F� �4^  Dу �`5  �� �� D-� �/M  �� �� 2)�A     �_  �]  3T1 2`�A     �_  �]  3T8 2ǁA     :^  ^  3Qq  G�A     '`  3T83Q	��B     3R
  �0  B� ���A     N       ��^  C.� �4^  ԭ Э C�  �
�  � 
� H� ��   QCV� ��   H� D� Dr� �
�   �� ~� D@�  �
�   � � Dm�  ��  � �  IEP  ��A     T       ��_  JWP  =� 5� KdP  KqP  LEP  �  JWP  �� �� M�  ?dP  � � ?qP  � � 2�A     �_  ^_  3Uv  7;�A     3`  3Us 3Tv 3Q8    N� � 	6N� � BN� � 	7	N��  ��  %7Nj j <O� � ( N�{ �{ =N� � GN��  ��  CN  &'	N�q  �q  J	N�} �} ?NaH aH %%	N��  ��  dN�� �� 	<	N� � ' �Q   ̩  S#  �� �*  ��A     =      �9 u�  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �  
K   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
K   /  ��   [r  �4 #�  �   �X  5�  
K   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K&  
�   P�  =_  ��   R�  N�  ��  ��   �p  W�  
K   3�  ��   ({  ��  ğ   F]  8�  
K   Y@  ��   �c  |  ��  l  ��  �   
K   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {@  
K   ��  &�   �  º  GY  �f  ��   v�  ��  
K   �  GQ   ϼ  �  �_  X  &�  �b   	"|  	*y  	��  	+y  	I�  	,y  	�a  	-y  
 	�  ��  
";   E�  
#;  e% 
$B  u  
%
�  �8 
&
�  ��  
)
�  /b  
-
�  ��  
.	�   a  
2
�  �T  
3
�   Mx 
4E  �  
K   ")  ��  WH  �~  �O  �m  ��   �  ��  ��  	 =� 5  ��  .j  ^�  2�   }�  7�  �� ;K    	�  r�  �   .� $�  O� )�   �  �  �    )  �  �  �   �  1   �  �  K   R   1    �  ��  ,j  �  �  oS  '  dS  ()k  � +
k   � ,�  @�  -
�   >z .
�   �  /R   �H  3{    �   {  =      	�� 7{  	�� 8K   t�   �   �  �  �  =   �' �  	��  1�  	]  4�  �  �  �  =   � �  	Zy  8�  �    =   =   �    	��  ;  Ʃ  QK   '  3  I  =     8  	�  WI  �p  #f  l  s   S�  $  �  �  R    T}  %�  �  �  R   R    '	�  acv )Z  ��  *s  ��  +�   �y -�  �Y  6�  ��  :-  s�  <-   �H  =-  xz  >�   �  x @�  B  O  =    4  _  =    
�	�  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x �_  
K     @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  
K   ��%  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u  (x	&   �u z    � {	�    s |	�    � ~�   N�  �%   ��  �	�    ��  �	�     J]  ��%  &  .&  =   � !�^  �&  �   F&  " !�  �;&  #K   ��)  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  S&  \	�*   �Y  	�     *O  	�    ��  	�    �  	�    b�  	�    ��  	�    �  	�    +�  	�    Zp  	�     o�   	�   $ m�  !	�   ( 4�  "	�   , �  #	�   0 �  $	�   4 ��  %	�   8 L� &	�   < ��  '	�   @   (	�   D ��  )	�   H \q *	�   L z�  +	�   P �  ,	�   T /�  -	�   X ʤ  /�)  �*  +  =   � !��  1+  �]  ���,  `e �3   x ��  y ��  z ��   ��  ��,  (cN  ��,  0Mp �'  8�u �  <� ��   @�H  ��,  Hr�  ��,  P��  �4-  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� ��)  �y� �:-  �s ��   ��� �@-  ��  ��   ��  ��   �ʺ  ��   ��l  ��   �  �  �,  � ��  �   � ��  	�   � �R   /  � f�  �   � I}  �  � ��  �,  � #+  Gx  �4-  >} ��2   �}  �B  �|  �B  
 �,  �*  &  $d  HN /  mo P�1   ��  Q�8  cmd R�  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g�8  8�W  h�8  P��  iy  h�� l�1  l�N  m�  |E�  p�  ��W  r�8  �~�  s�1  �*� t�1  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��1  �%�R  ��    %��  ��   %�  ��   %h  ��8  %I�  �y  @ F-  �z #+  	��  ��   	�\  �y  	�  �W/  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  ��  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   (	90  ��  B      B  Vd  !B  �  "B  �� #90   �   I0  =    � %�/  C	u0  x E�   y F�   �{ HU0  (T	�0  `e V3   x W�  y X�  z Y�    	�  [�0  �a	�1  = c�   F�  d�  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  o�1  ��  r
�1   iK  u�0  0��  x
�   XS�  {�1  `��  ~R   h��  ��   pu| �u2  x &/  �   �1  =    �}  X�u2  v1 �*3   v2 �*3  dx ��  dy ��  �  �B  �k �B  tag �B  �W  �?  �o �03  $��  �3  4SX  ��2  8d�  ��2  @��  �
�   H��  �R   P {2  �1  �z ��0  �	�2  2�  ��   ]  ��  �h  �B  �N  �B  
�K  �B  >} ��2   �2  �}  ��2  
K   �3  ��   �  o�  ��   ��  ��2  u0  �  @3  =    �u  ��1  �z ��,  8�	�3  v1 �*3   v2 �*3  82  ��  Mp �'  [�  ��3   �  ��3   SX  ��2  (d�  ��2  0 �2  @3  A{ �X3  4	94  &x �   &y 	�  &dx 
�  &dy �   �o 94   )�  O  0 �  O4  =   =    (} �3  �  *�  'v  @25   @�  45   &x1 5�   &x2 6�    .]  8�   5]  9�   �� :�   ��  =�    �  @�    ��  C�  $ �n  G$5  ( 9x  H$5  0 �^  I$5  8 �3  B  >�  Ki4  '�h  PR6   s�  U6    �H  V6  &x1 X�   &x2 Y�   &gx \�  &gy ]�  &gz `�   &gzt a�  $ �x  d�  ( � f�  , ~�  i�  0 t  k�  4 .� l�   8 �  p6  @ 	�  r�   H 75  \4  �h  t75  �	a6   �c  �y    �O  �a6   �x  �
q6   B  q6  =    �  �6  =    I�  �,6  �	�6   �  ��     �  ��6   �6  �  ��6  (��	r7     ��    �  �	�    t�  �	�    ��  �	�    /�  �	�    �  �	�  &top �	r7  )��  �	�  U)��  �	�  V)� �	r7  W)�  �	�  � �  �7  =   ? ��  ��6  	�7  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�7  �7  8  =    	S�  '�7  
K   718  {�   U�  ~�   >	m8  �� @@-   s A
�   sx B�  sy C�   Nz E18  
K   1�8  ��   ��  ��   �y  9y8  �   �8  =    y  �8  =    y  �8  =    m8  �8  =    hy �F-  (�	V9  in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�1  �a  �
�   $ ��  ��8  ��	�9  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��9  ( V9  :  =    ޴  �b9  	.L  &#:  �  	׮  )#:  	�  +#:  	�  ,#:  	�Q  .6  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�:  �   	��  8�:  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�:  �6  	��  H�   	��  I*3  	��  K�   	a� L5  	w�  N�   	P{ O�2  	��  Q�   	��  RI;  L3  	��  T�   	�� Ug;  O4  	�}  W�   	u| X�3  	M�  Z�   	P�  [�3  	��  a�  	��  b�  	�  c�  	�p  e'  	�T  f�;  �8  	�a  j'  �   �;  =   � 	ը  l�;  '  <  =   @ 	�p  m<  	 �  p�  	p|  q'  	$Y  v�   	�K  y�   	g  {a<  �7  	d�  |a<  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   6  =  =   =   / 	��  E=  6  5=  =   / 	Ԁ  F%=  6  W=  =   =    	7� GA=  	�R  I�   	��  J6  	��  U�   	P�  \�  	��  ]�  	L�  ^�  	ߵ  _�  	�  a�  	@�  5  	[�  �3  	 �  �3  	SX  �2  	d�  �2  	��  �   	_�   �   	��  "y  	��  %y  	'�  &y  	�]  (y  *5  W>  =   � 	�P  *G>  	ӯ  +o>  *5  	|  -�>  6  	��  .�>  	��  /�>  �>  �>  �   �    	��  $5  �   �>  	qY  "�>  	�  #�>  B  �>  =   ? 	��  %�>  	��  &�>  �  ?  =   � 	@Y  (?  �  ;?  =   ? 	V�  )*?  6  W?  =    	�h  G?  	�  o?  6  	�  6  	�f  !�>  	r�  "�>  	��  %$5  	��  &$5  	׆  '�  	��  (�  	�  *�  	��  +�  	�  6  	��  �   	�_  �   	�_  �   	b  �  	t  �  	j�  "�  	�  :�   	��  ;�   	��  <�   	�W  >6  	hn  @�  	U~  A�  	�  B�  	 �  C�  	%�  F�  	�u  H�  	z  I�  	N�   %�1  	��   '�  I0  �  	��  !My  	(h  !N�   	l�  !N�   	�  ".y  	�  "/y  	�  "0y  	�  "2y  	w�  "8  	�  "9�  	�  ":�  	�_  ";�   	��  ">y  	�  "Jy  	"�  "R�  	t�  "S�   	�w  "T�   	؜  "Y�   	q�  "[y  	Ƚ  "^�  	�  "_�   	�y  "`�   	b�  "c�   	+�  "fy  	��  "iy  	֘ "l�   	�J  "x�   	��  "y�   	ks  "�   	�  "��   	J�  "��   	�i  "��   	��  "�y  	��  "�y  	��  "�y  	<� "�y  	��  "�y  	��  "�y  	5�  "�y  	<m  "��   	 K  "��   	�R  "��   	op  "��   	�m  "��   	D  "��   	X�  "��   	If  "��   	� "��   	��  "�y  	�U  "�y  	`  "�y  	J�  "�y  	��  "�y  	� "��  �8  iC  =    	�  "�YC  y  �C  =    	� "�uC  �  �C  =   	 	,�  "��C  	R�  "��C  �  �  �C  =    	�u  "��C  	��  "�:  	�e  "��   �   D  =   � 	(�  "��C  	�  "�y  !��  "�  !�v  "�   !n�  "�   !4�  "�   !*b "�   !��  "�@  *� 9�  	h�f     +Y:  :	��f     +e:  ;	@�f     +q:  <	X�f     +�<  =	`�f     +�<  >	D�f     �  �D  =   ? *h� ?�D  	`�f     �   E  =   _ *�� @E  	��f     �  >E  =   =   � *�� F(E  	��f     ,� K�  	��e     +�?  R	��f     +�?  S	��f     +�?  T	��f     +@  U	��f     +@  V	p�f     +@  W	H�f     +)@  Z		��f     *p� ]�   	��f     �   F  =   1 -�� �E  	`be     --� �   	��e     .�@  �	��f     .�@  �	��f     .5@  :	x�f     .A@  ;	|�f     .M@  <	t�f     .Y@  >	��f     .e@  @	L�f     .q@  A	��f     .}@  B	��f     .�@  C	��f     .�@  F		P�f     -Z� I�   	d�f     /Y ���A     �       �H  0top �
�   _� [� 1<p �
�   �� �� 0ofs �
�   հ ϰ 0i �
�   5� 3� 2ИA     H  �G  3U03T{  2�A     H  �G  3T{  2�A     H  �G  3Ux 3Ty  41�A     2Q  3U03T03Q
@3R�  /�1 �`�A     %       �XH  5ofs �K   \� X� 6r� ��   �� ��  /� ,�A     q      �7K  0src .�  � � 1`5 /�  � � 0x 0
�   �� �� 0y 1
�   =� /� 1.� 2�@  � ׳ 7F� 5�   
T�B     �7L� 8�   
L�B     �1� :�   �� �� 8�A     >Q  29�A     JQ  QI  3U
 �3T13Q0 2_�A     VQ  hI  3T8 8��A     bQ  2ǖA     VQ  �I  3U	]�B     3T8 2�A     nQ  �I  3Qv  2�A     VQ  �I  3U	d�B     3T8 2+�A     nQ  �I  3Qv  2>�A     VQ  J  3U	k�B     3T8 2e�A     nQ  )J  3Qv  2x�A     VQ  MJ  3U	r�B     3T8 2��A     nQ  eJ  3Qv  2��A     VQ  �J  3U	y�B     3T8 8͗A     nQ  2ܗA     VQ  �J  3U	��B     3T8 8��A     nQ  2�A     VQ  �J  3U	��B     3T8 8%�A     nQ  24�A     VQ  K  3U	��B     3T8 8T�A     nQ  9\�A     zQ   /ƅ 	��A     f       ��K  :��  
�   U:  �   T0i 
�   �� ��  /� ���A           �VL  1@�  �K   J� F� 1r� �K   �� �� 1b� �K   �� �� 1�� �K   � � 1`5 ��  +� %� 1r� �	�   |� v� 1�q �	�   ɶ Ƕ ;A     �Q  3U	1�B       /�� N��A     �       �$M  1@�  PK   �� �� 1r� PK   5� 3� 1`5 Q�  Z� X� 1r� R	�   �� }� 1�q S	�   з η 1b� TK   �  � 1�� TK   B� >� ;�A     �Q  3U	1�B       /҆ �A     �       �vM  0i 
�   �� �� ;/�A     JQ  3U
 3T13Q0  /�� �#�A     �       �3N  1r� ��   ޸ ָ 1`5 ��  I� A� 1M9 ��  �� �� 1{q ��  3� -� 1n� ��  ~� |� 0x ��   �� �� ;m�A     �Q  3U	��B     3Rs   /C� �h�A     �       ��N  1r� ��   � ݺ 1`5 ��  N� H� 1{q ��  �� �� 1n� ��  � � ;��A     �Q  3U	��B       /�� VO�A           �qO  1r� X�   � � 1`5 Y�  � y� 1M9 Z�  Ѽ ˼ <{q [�  1n� \�  � � 0x ]	�   N� J� ;ƐA     �Q  3U	�B       /x� v�A     �       ��O  1r� �   �� �� 1`5 �  �� � <{q �  1n�  �  E� C� ;�A     �Q  3U	�B       =�� ���A     �       ��P  >r� ��   x� p� >`5 ��  � ۾ >M9 ��  Y� Q� >{q ��  Ϳ ǿ >n� ��  � � ?x ��   A� ;� ;�A     �Q  3U	��B       =� f��A     �       �2Q  >r� h�   �� �� >`5 i�  
� � >{q j�  \� V� >n� k�  �� �� ;:�A     �Q  3U	��B       @��  ��   E@� � 7	@� � 6@��  ��  C@w� w�  R@y�  y�   9@� �  V@��  ��  #7 wJ   s�  S#  �� �*  2�A     J	      II =�  �)  �=   ,	  int ^&  9�  �� �  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2D   8;:  5D   < �   1  �K 8"p   	�  K     	�  L  	�  M  0t  B  e2    �0  }  ��  6  
i   J�  D   �C  
D  ���� �C  Nj  ڵ  R^  �  
i   Y�  ��   �c  |  ��  l  ��  �   
i   k5  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {�  
i   �t  &�   �  º  GY  �f  ��   v�  �A  
i   ��  GQ   ϼ  �  �_  X  &�  �b    	E  ��  "P   E�  #P  e% $W  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	D   a  2
�  �T  3
�   Mx 4�  �  ^   W  	��  	M�  	(h  	ND   	l�  	ND   t�  
 D   �  
i   �  �L  M M �L  	B 8D   	x	 9D   �  �  =   �' �  	��  1�  	]  4  �  �    =   �   	Zy  8  �  D  =   =   � .  	��  ;D  Ʃ  Qi   U  a  w  =     f  	�  Ww  �p  #^  S�  $�  �  �  K    T}  %�  �  �  K   K    '	  acv )�  ��  *�  ��  +�   �y -�  �Y  6  ��  :N  s�  <N   �H  =N  xz  >     x @  W  p  =    I  �  =    
�	�  x �W   y �W  Mp �W  *� �W  ޽  �W   ~x ��  
i   $	  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  
i   ��"  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u0	  (x	1#  �u z$	   � {	D   s |	D   � ~  N�  �"  ��  �	D   ��  �	D     J]  ��"  1#  O#  =   � �^  �>#  �   g#   �  �\#   i   ��&  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  t#  \	(  �Y  	D    *O  	D   ��  	D   �  	D   b�  	D   ��  	D   �  	D   +�  	D   Zp  	D    o�   	D   $m�  !	D   (4�  "	D   ,�  #	D   0�  $	D   4��  %	D   8L� &	D   <��  '	D   @  (	D   D��  )	D   H\q *	D   Lz�  +	D   P�  ,	D   T/�  -	D   X ʤ  /�&  (  7(  =   � ��  1'(  �]  ��*  `e �T   x ��  y ��  z ��   ��  �*  (cN  �*  0Mp �U  8�u �$	  <� �D   @�H  �*  Hr�  �*  P��  �U*  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  �D   |*� ��&  �y� �[*  �s �D   ��� �a*  ��  �D   ��  �D   �ʺ  �D   ��l  �D   � �  *  ���  D   ���  	D   ��R  A,  �f�  D   �I}  �  ���  *  � D(  Gx  �U*  >} ��/   �}  �W  �|  �W  
  *  (  1#  !d  HNA,  mo PR.   ��  QM5  cmd RE  �  W�  (_  Y�   #_  [�  $bob ]�  (�  aD   ,�[  bD   0sb  dD   4d]  gY5  8�W  hi5  P��  i�  h�� lX.  l�N  m5  |E�  p5  ��W  ry5  �~�  sX.  �*� tX.  ��� wD   ���  xD   �X�  |D   ��e  D   ���  �D   �g  �D   ��u  �D   �|G ��   �Q  �D   ��  �D   �o�  �R.  �"�R  �D    "��  �D   "�  �D   "h  ��5  "I�  ��  @ g*  �z D(  	��  ��   	�\  ��  	�  �b   	��  �D   	��  �D   	2�  ��  	��  �D   	Ɇ  �Q  	��  �D   	��  �D   	�h  �D   	rK  �D   	l�  �D   	]�  �D   	��  �D   C	(-  x E�   y F�   �{ H-  (T	l-  `e VT   x W�  y X�  z Y�    	�  [4-  �a	R.  = c�   F�  d�  �~ eW  h�  fW  
t�  gW  �k hW  tag iW  �N  l
D   ��  oR.  ��  r
X.   iK  ul-  0��  x
D   XS�  {R.  `��  ~K   h��  �D   pu| �(/  x G,  D   h.  =    �}  X�(/  v1 ��/   v2 ��/  dx ��  dy ��  �  �W  �k �W  tag �W  �W  �`  �o ��/  $��  ��/  4SX  ��/  8d�  ��/  @��  �
D   H��  �K   P ./  h.  �z �x-  �	�/  2�  ��   ]  ��  �h  �W  �N  �W  
�K  �W  >} ��/   4/  �}  �@/  
i   ��/  ��   �  o�  ��   ��  ��/  (-  �  �/  =    �u  �h.  �z � *  8�	{0  v1 ��/   v2 ��/  82  ��  Mp �U  [�  �{0   �  ��0   SX  ��/  (d�  ��/  0 �/  �/  A{ �0  4	�0  #x �   #y 	�  #dx 
�  #dy �  �o �0  )�  p  0 �  1  =   =    (} �0  �  *�  $v  @2�1  @�  4�1   #x1 5D   #x2 6D   .]  8�  5]  9�  �� :�  ��  =D   �  @�   ��  C�  $�n  G�1  (9x  H�1  0�^  I�1  8 �0  W  >�  K1  $�h  PR�2  s�  U�2   �H  V�2  #x1 XD   #x2 YD   #gx \�  #gy ]�  #gz `�   #gzt a�  $�x  d�  (� f�  ,~�  i�  0t  k�  4.� lD   8�  p�2  @	�  rD   H �1  1  �h  t�1  �	3  �c  ��   �O  �3  �x  �
$3   W  $3  =    �  43  =    I�  ��2  �	h3  �  �D    �  �h3   43  �  �A3  %��	%4    ��   �  �	D   t�  �	D   ��  �	D   /�  �	D   �  �	�  #top �	%4  &��  �	�  U&��  �	�  V&� �	%4  W&�  �	�  � �  64  =   ? ��  �{3  	�4  ~�  t   �S  
D   ��   
D     !
D   �g  "
D   �^  #
D    ��  %C4  �4  �4  =    	S�  '�4  
i   7�4  {�   U�  ~�   >	 5  �� @a*   s A
D   sx B�  sy C�   Nz E�4  
i   1M5  ��   ��  ��   �y  9,5  D   i5  =    �  y5  =    �  �5  =     5  �5  =    hy �g*  	.L  &�5  �  	׮  )�5  	�  +�5  	�  ,�5  	�Q  .�2  	��  0D   	��  1D   	(_  2D   	դ  4D   	�j  7#6  D   	��  8#6  	@�  <D   	�O  =D   	(g  >D   	�^  ED   	�u Fq6  n3  	��  HD   	��  I�/  	��  KD   	a� L�1  	w�  ND   	P{ O�/  	��  QD   	��  R�6  �/  	��  TD   	�� U�6  1  	�}  WD   	u| X�0  	M�  ZD   	P�  [{0  	��  a�  	��  b�  	�  c�  	�p  eU  	�T  fg7  �5  	�a  jU  D   �7  =   � 	ը  ly7  U  �7  =   @ 	�p  m�7  	 �  p�  	p|  qU  	$Y  vD   	�K  yD   	g  {�7  64  	d�  |�7  	��   �  		�  !�  	�3 #D   	_  $D   	-�  (D   	�f  )D   	�G  +�  	`�  ,�  	A�  -�  	��  /D   	��  1D   	P�  2D   �2  �8  =   =   / 	��  E�8  �2  �8  =   / 	Ԁ  F�8  �2  �8  =   =    	7� G�8  	�R  ID   	��  J�2  	��  UD   '	P�  \"9  9  	��  ]"9  	L�  ^"9  	ߵ  _"9  	�  a"9  	@�  �1  	[�  {0  	 �  �0  	SX  �/  	d�  �/  	��  D   	_�   D   	��  "�  	��  %�  	'�  &�  	�]  (�  �1  �9  =   � 	�P  *�9  	ӯ  +:  �1  	|  -:  �2  	��  .:  	��  /:  ::  J:  D   D    	��  �1  �   4:  	qY  "V:  	�  #V:  W  �:  =   ? 	��  %z:  	��  &z:  �  �:  =   � 	@Y  (�:  �  �:  =   ? 	V�  )�:  �2  �:  =    	�h  �:  	�  ;  �2  	�  �2  	�f  !z:  	r�  "z:  	��  %�1  	��  &�1  	׆  '�  	��  (�  	�  *�  	��  +�  	�  �2  	��  D   	�_  D   	�_  D   	b  �  	t  �  	j�  "Q  	�  :D   	��  ;D   	��  <D   	�W  >�2  	hn  @�  	U~  A�  	�  B�  	 �  C�  	%�  FQ  	�u  HQ  	z  IQ  	- D   	_   D   ( K  /D   	zg     )m8  2	(ce     )�8  5	 zg     	� 6:  )18  8	@g     )=8  9	�f     )I8  ;	��f     )U8  <	��f     )a8  =	�f     (y� @D   	��f     )�7  B	��f     )y8  C	�4g     )�8  D	��f     )+7  F	zg     )77  G	zg     )C7  H	zg     )O7  J	�f     )8  L	�f     )8  M	��f     )[7  O	�4g     )	9  R	��f     )m7  W	�f     )�7  ]	@�f     )�7  b	 ug     )�8  d	�g     )�8  e	`g     )�8  f	 5g     )�8  i	��f     )9  m	��f     )49  n	zg     )@9  o	 �f     )(9  p	��f     )L9  q	 �f     *� �
�  	��f     *`� �D   	zg     *4� �D   	��f     +� _5�A     G       ��?  ,�R  _$g7  �� �� -;�A     �?  K?  .Uu  /@�A     �I  /E�A     �I  /J�A     �I  /O�A     �I  /T�A     �I  /b�A     �I  /g�A     �I  /l�A     �I  /q�A     �I  /v�A     J  0|�A     �I   +Z� 7v�A     �       �@  1�R  7g7  U2i 9
D   � �  33, �6  �A     ]       ��@  4x �  I� C� 4y �  �� �� 5=� �6  �� �� 5<p 
D   � � 5	�  
D   5� 1� 6X�A     _H  .Uv .T| .Qs   +C ���A     �       ��A  7�B  ��A     ��A     "       	A  8�B  8�B   /��A     J  -��A     J  ;A  .U. -��A     J  SA  .U. -��A     J  kA  .U. /�A     &J  -�A     J  �A  .U. /�A     �B  -��A     J  �A  .U. /��A     2J  /�A     >J  6�A     J  .U.  +�	 ��A     �      ��B  9� ��  2dy ��  o� k� 2i �
D   �� �� 2j �
D   �� |� 5� �
D   �� �� 5�w  �
D   e� a� /C�A     JJ  /H�A     |C  /ϟA     VJ  6�A     VJ  .U@<$  :�[ ��B  ;=g �D   ;��  �D    +.� bu�A     �       �|C  2i d
D   �� �� 2j e
D   �� �� 5� f
D   � � 5�w  g
D   �� �� 5� h
D   �� �� 6��A     VJ  .UDC$.Tv D$  +K� f�A           �#D  2i D   3� 1� 2x D   ^� V� 2t  D   �� �� 5m� !�  [� W� /��A     VJ  -��A     bJ  D  .Ts  6-�A     bJ  .Ts   <!� �3�� �	�  ݛA     �       �"E  ,� �)U  �� �� 5� ��  �� �� 5@� �U  �� �� 9� �U  5�� �D   T� R� 9g� �D   2num ��  {� w� 2den �D   �� �� /�A     bJ  --�A     bJ  E  .Ts  6D�A     VJ  .Uv   <G� �3� x�  w�A     e       ��E  4x y�  �� �� 4y z�  D� @� 9Mp |
D   2dx }�  �� }� 2dy ~�  �� �� 9v� �  9S� ��  5{q ��  Q� M� -��A     VJ  �E  .Ts  0ܛA     VJ   3Ef jU  b�A            ��F  4x1 k�  �� �� 4y1 l�  �� �� 4x2 m�  ?� ;� 4y2 n�  |� x� =w�A     �F  .U�Q.T�R  3w� U  W�A           �AG  4x �  �� �� 4y �  �� �� /��A     nJ  /��A     nJ  /ȚA     nJ  /ߚA     nJ  /�A     nJ  /�A     nJ  /9�A     nJ  /P�A     nJ   >ɇ �D   әA     �       �_H  ?x ��  �� �� ?y ��  :� 4� @��  �
�1  �� �� Alx ��  �� �� Aly ��  � �� Aldx ��  G� 7� Aldy ��  � 
� Adx ��  H� D� Ady ��  �� ~� BϷ  ��  �� �� B�T  ��  	� � /<�A     bJ  6H�A     bJ  .Uv .Ts   >� �D   Q�A     �       �)I  ?x ��  2� ,� ?y ��  �� ~� @=� ��6  �� �� Adx ��  9� 7� Ady ��  `� \� BϷ  ��  �� �� B�T  ��  �� �� /��A     bJ  6ęA     bJ  .Uv   C�� {2�A            �nI  Dx |D   UDy }D   TDbox ~�5  Q E"E  ܛA            �F�B  ��A            ��I  G�B  UG�B  T H� � 6H� � 7H� � ,H�� �� 7H��  ��  	7Hf� f� :H� � <H>� >� 8Hƃ ƃ $I� �  H�� �� +H'� '� #H҆ ҆ \Hƅ ƅ UHH_  H_  
#	Hd  d  
"	H�� �� \ 2K   ܱ  S#  u� �*  |�A           UW ��  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  9�  0t  4  e2    �0  }  ��  (  
K   J�  D   �C  
D  ���� �C  N\  ڵ  RP  �   	)  ��  "B   E�  #B  e% $I  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�  ;  
K   "�  ��  WH  �~  �O  �m  ��   �  ��  ��  	 
K   	�  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  	(�  
K   	/  ��   [r  �4 #�  �   �X  	5�  
K   	:t  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  	K  
�   	P�  =_  ��   R�  N�  ��  ��   �p  	W�  =� 
�  ��  
.   ^�  
2�   }�  
7�  �� 
;K    
	1  r� 
 F   .� 
$W  O� 
){   @  @  �    �  1  W  @   L  1   {  @  K   R   1    ]  ��  
,   �  �  oS  '�  dS  ()  � +
   � ,@  @�  -
�   >z .
�   �  /R   �H  3    �     =    �  	�� 7  	�� 8K   
K   3V  ��   ({  ��  ğ   F]  8/  
K   Y�  ��   �c  |  ��  l  ��  �   
K   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {�  
K   �+  &�   �  º  GY  �f  ��   v�  ��  
K   �p  GQ   ϼ  �  �_  X  &�  �b   I  �  =    ;  �  =    
�	�  x �I   y �I  Mp �I  *� �I  ޽  �I   ~x ��  �   �  )  	��  M�  	(h  N�   	l�  N�   	r  ~�  +   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %  r  �  =    	S�  '~  t�   �   �  �  �  =   �' �  	��  1�  	]  4�  �  �  �  =   � �  	Zy  8�  �    =   =   �   	��  ;  Ʃ  QK   (  4  J  =     9  	�  WJ  �p  #�  S�  $s  y  �  R    T}  %�  �  �  R   R    '	�  acv )[  ��  *g  ��  +�   �y -�  �Y  6�  ��  :!	  s�  <!	   �H  =!	  xz  >�   �  x @�  
K   �  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �3	  
K   �&  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�  (x	�&   �u z�    � {	�    s |	�    � ~�   N�  &   ��  �	�    ��  �	�     J]  �$&  �&  �&  =   � !�^  ��&  �   �&  " !�  ��&  #K   � *  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �&  \	z+   �Y  	�     *O  	�    ��  	�    �  	�    b�  	�    ��  	�    �  	�    +�  	�    Zp  	�     o�   	�   $ m�  !	�   ( 4�  "	�   , �  #	�   0 �  $	�   4 ��  %	�   8 L� &	�   < ��  '	�   @   (	�   D ��  )	�   H \q *	�   L z�  +	�   P �  ,	�   T /�  -	�   X ʤ  /-*  z+  �+  =   � !��  1�+  
K   7�+  {�   U�  ~�   >	,  �� @,   s A
�   sx B�  sy C�   �&  Nz E�+  �]  ���-  `e �'	   x ��  y ��  z ��   ��  ��-  (cN  ��-  0Mp �(  8�u ��  <� ��   @�H  ��-  Hr�  ��-  P��  �$.  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� � *  �y� �*.  �s ��   ��� �,  ��  ��   ��  ��   �ʺ  ��   ��l  ��   �  �  �-  � ��  �   � ��  	�   � �R  
0  � f�  �   � I}  �  � ��  �-  � ,  Gx  �$.  >} �o8   �}  �I  �|  �I  
 �-  z+  $d  HN
0  mo PJ0   ��  Q>0  cmd R)  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  gP0  8�W  h`0  P��  i�  h�� lp0  l�N  m�  |E�  p�  ��W  r�0  �~�  sp0  �*� tp0  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �J0  �%�R  ��    %��  ��   %�  ��   %h  ��0  %I�  ��  @ 0.  �z ,  
K   1>0  ��   ��  ��   �y  90  0  �   `0  =    �  p0  =    �   �0  =    �  �0  =    ,  �0  =    hy �0.  (�	1  in ��   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
p0  �a  �
�   $ ��  ��0  ��	�1  2�  �
�    I�  ��  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��1  ( 1  �1  =    ޴  �1  	�  .�  	�  /�  	�  0�  	�  2�  	w�  8  	�  9�  	�  :t  	�_  ;�   	��  >�  	�  J�  	"�  R�  	t�  S�   	�w  T�   	؜  Y�   	q�  [�  	Ƚ  ^�  	�  _�   	�y  `�   	b�  c�   	+�  f�  	��  i�  	֘ l�   	�J  x�   	��  y�   	ks  �   	�  ��   	J�  ��   	�i  ��   	��  ��  	��  ��  	��  ��  	<� ��  	��  ��  	��  ��  	5�  ��  	<m  ��   	 K  ��   	�R  ��   	op  ��   	�m  ��   	D  ��   	X�  ��   	If  ��   	� ��   	��  ��  	�U  ��  	`  ��  	J�  ��  	��  ��  	� �V  �0  94  =    	�  �)4  �  U4  =    	� �E4  �  q4  =   	 	,�  �a4  	R�  ��4  �  �  �4  =    	�u  ��4  	��  ��1  	�e  ��   �   �4  =   � 	(�  ��4  	�  ��  !��  V  !�v  �   !n�  �   !4�  �   !*b �   !��  �  	��  ��   	�\  ��  	�  �^5  �  	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  ��  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	6  x E�   y F�   �{ H�5  (T	Y6  `e V'	   x W�  y X�  z Y�    	�  [!6  �a	?7  = c�   F�  d�  �~ eI  h�  fI  
t�  gI  �k hI  tag iI  �N  l
�   ��  oJ0  ��  r
p0   iK  uY6  0��  x
�   XS�  {J0  `��  ~R   h��  ��   pu| ��7  x �}  X��7  v1 ��8   v2 ��8  dx ��  dy ��  �  �I  �k �I  tag �I  �W  �p  �o ��8  $��  ��8  4SX  �o8  8d�  �o8  @��  �
�   H��  �R   P 8  ?7  �z �e6  �	o8  2�  ��   ]  ��  �h  �I  �N  �I  
�K  �I  >} �o8   8  �}  �8  
K   ��8  ��   �  o�  ��   ��  ��8  6  �  �8  =    �u  �?7  �z ��-  8�	R9  v1 ��8   v2 ��8  82  ��  Mp �(  [�  �R9   �  �X9   SX  �o8  (d�  �o8  0 u8  �8  A{ ��8  4	�9  &x �   &y 	�  &dx 
�  &dy �   �o �9   )�  �  0 �  �9  =   =    (} j9  �  *�  'v  @2�:   @�  4�:   &x1 5�   &x2 6�    .]  8�   5]  9�   �� :�   ��  =�    �  @�    ��  C�  $ �n  G�:  ( 9x  H�:  0 �^  I�:  8 ^9  I  >�  K�9  '�h  PR�;   s�  U�;    �H  V�;  &x1 X�   &x2 Y�   &gx \�  &gy ]�  &gz `�   &gzt a�  $ �x  d�  ( � f�  , ~�  i�  0 t  k�  4 .� l�   8 �  p�;  @ 	�  r�   H �:  �9  �h  t�:  �	�;   �c  ��    �O  ��;   �x  �
�;   I  �;  =    �  <  =    I�  ��;  �	?<   �  ��     �  �?<   <  �  �<  (��	�<     ��    �  �	�    t�  �	�    ��  �	�    /�  �	�    �  �	�  &top �	�<  )��  �	�  U)��  �	�  V)� �	�<  W)�  �	�  � �  =  =   ? ��  �R<  	.L  &&=  �  	׮  )&=  	�  +&=  	�  ,&=  	�Q  .�;  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�=  �   	��  8�=  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�=  E<  	��  H�   	��  I�8  	��  K�   	a� L�:  	w�  N�   	P{ Oo8  	��  Q�   	��  RL>  �8  	��  T�   	�� Uj>  �9  	�}  W�   	u| XX9  	M�  Z�   	P�  [R9  	��  a�  	��  b�  	�  c�  	�p  e(  	�T  f�>  �0  	�a  j(  �   �>  =   � 	ը  l�>  (  ?  =   @ 	�p  m?  	 �  p�  	p|  q(  	$Y  v�   	�K  y�   	g  {d?  =  	d�  |d?  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   �;  @  =   =   / 	��  E@  �;  8@  =   / 	Ԁ  F(@  �;  Z@  =   =    	7� GD@  	�R  I�   	��  J�;  	��  U�   	P�  \5  	��  ]5  	L�  ^5  	ߵ  _5  	�  a5  	@�  �:  	[�  R9  	 �  X9  	SX  o8  	d�  o8  	��  �   	_�   �   	��  "�  	��  %�  	'�  &�  	�]  (�  �:  ZA  =   � 	�P  *JA  	ӯ  +rA  �:  	|  -�A  �;  	��  .�A  	��  /�A  �A  �A  �   �    	��  �:  �   �A  	qY  "�A  	�  #�A  I  �A  =   ? 	��  %�A  	��  &�A  �  !B  =   � 	@Y  (B  �  >B  =   ? 	V�  )-B  �;  ZB  =    	�h  JB  	�  rB  �;  	�  �;  	�f  !�A  	r�  "�A  	��  %�:  	��  &�:  	׆  '�  	��  (�  	�  *�  	��  +�  	�  �;  	��  �   	�_  �   	�_  �   	b  �  	t  �  	j�  "�  	�  :�   	��  ;�   	��  <�   	�W  >�;  	hn  @�  	U~  A�  	�  B�  	 �  C�  	%�  F�  	�u  H�  	z  I�  	-  �   	_    �   *�A  %	X�h     +ӈ &�A  	P�h     =  D  =    +�� .�C  	 �g     +>� /d?  	H�h     *X?  0	`�h     *j?  1	��g     I  mD  =   �O +ʈ 5	\D  	��h     *�A  6
	 �g     *�A  >		��g     *B  ?		��i     �   �D  =   � +�� E�D  	 �g     +�� F�D  	`}g     +2� K�A  	��g     +�� L�  	@�g     *!B  N	 �h     *>B  O	 �g     +߈ P�  	 �g     +�� Q�  	@�h     +h� SB  	��g     +v� TB  	@zg     +&� UB  	��g     +\� VB  	`�g     ,� ho�A           �G  -pl jd?  �� �� .�R  k�   � � -x l�   p� f� .�� m�   �� �� .Mp n�   � � .C� o�   -� +� /��A     �J  �F  0U	��B      /ӦA     �J  �F  0U	��B      /��A     �J  �F  0U	�B      1��A     �J  /ͧA     K  �F  0Uv 0T1 1e�A     G  2n�A     K  0Uv   3j� D��A     �       ��G  4x E�   V� P� 4t1 F�   �� �� 4b1 G�   @� 4� 4t2 H�   �� �� 4b2 I�   G� =� /�A     tI  �G  0U 0Q��� 2)�A     tI  0Q}   5�� d?  =�A            ��H  4pl d?  �� �� 6' �   T7�� �   <� 4� .K� 
�   �� �� .� 	
�   �� �� .�� 

�   �� �� .�� 
�   � � -x 
�   4� 0�  8M� �d?  ��A     �       �I  9  ��  n� j� 9�  ��   �� �� 9t�  ��   �� �� :Wy �d?  6� 0� 2��A     �J  0U	��B       ;� ��A     �       �tI  <i �
�   �� �� :Mp �(  �� �� 1��A     K  1��A     K   =Q� r}�A     �      ��J  >y s�   � � >x1 t�   l� f� >x2 u�   �� �� :Mp w(  � 
� :#�  x�  9� /� :�� y�  �� �� :�8 zK   �� �� /��A     �J  KJ  0U	��B     0Tv 0Q| 0R}  1�A     )K  /��A     )K  pJ  0Us  /�A     )K  �J  0Us  /Y�A     )K  �J  0Us  /��A     )K  �J  0T��� 2��A     )K  0T���  ?�� ^|�A            �@��  ��  !7@�� �� "@� � B@} } I	@H_  H_  #	@d  d  "	 I   ǵ  S#  �� �*  ��A     �      �` Ѭ  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  9�  0t  4  e2    �0  }  ��  (  
K   J�  D   �C  
D  ���� �C  N\  ڵ  RP  �   	)  ��  "B   E�  #B  e% $I  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�  ;  
K   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (<  
K   /�  ��   [r  �4 #�  �   �X  5�  
K   :/  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K�  
�   Pn  =_  ��   R�  N�  ��  ��   �p  W;  
K   	3�  ��   ({  ��  ğ   F]  	8z  
K   	Y�  ��   �c  |  ��  l  ��  �   
K   	k7  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  	{�  
K   	�v  &�   �  º  GY  �f  ��   v�  	�C  
K   	��  GQ   ϼ  �  �_  X  &�  �b   I  �  =    ;  �  =    

�	"  x 
�I   y 
�I  Mp 
�I  *� 
�I  ޽  
�I   ~x 
��  �  ;   4  )  	��  M�  	(h  N�   	l�  N�   	�  ~�  v   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %k  �  �  =    	S�  '�  t�   �   �  �    =   �' �  	��  1  	]  4*  �  �  A  =   � 0  	Zy  8A  �  h  =   =   � R  	��  ;h  Ʃ  QK   y  �  �  =     �  	�  W�  �p  #;  S�  $�  �  �  R    T}  %�  �  �  R   R    '	%  acv )�  ��  *�  ��  +�   �y -�  �Y  6%  ��  :r  s�  <r   �H  =r  xz  >1   =  x @=  
K   �
  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  
K   �h$  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�
  (x	�$  �u z�
   � {	�   s |	�   � ~%  N�  h$  ��  �	�   ��  �	�     J]  �u$  �$   %  =   �  �^  ��$  �   %  !  �  �%  "K   �q(  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  %%  \	�)  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /~(  �)  �)  =   �  ��  1�)  
K   7*  {�   U�  ~�   >	R*  �� @R*   s A
�   sx B�  sy C�   �$  Nz E*  �]  ��:,  `e �x   x ��  y ��  z ��   ��  �:,  (cN  �:,  0Mp �y  8�u ��
  <� ��   @�H  �:,  Hr�  �:,  P��  �u,  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� �q(  �y� �{,  �s ��   ��� �R*  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  :,  ���  �   ���  	�   ��R  [.  �f�  �   �I}  "  ���  :,  � d*  Gx  �u,  >} ��6   �}  �I  �|  �I  
 @,  �)  #d  HN[.  mo P�.   ��  Q�.  cmd R)  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g�.  8�W  h�.  P��  i�  h�� l�.  l�N  m7  |E�  p7  ��W  r�.  �~�  s�.  �*� t�.  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��.  �$�R  ��    $��  ��   $�  ��   $h  ��.  $I�  ��  @ �,  �z d*  
K   1�.  ��   ��  ��   �y  9n.  a.  �   �.  =    �  �.  =    �   �.  =    �  �.  =    X*  �.  =    hy ��,  (�	a/  in ��   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�.  �a  �
�   $ ��  ��.  ��	0  2�  �
�    I�  ��  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  �0  ( a/  0  =    ޴  �m/  	�  .�  	�  /�  	�  0�  	�  2�  	w�  8�  	�  9�  	�  :/  	�_  ;�   	��  >�  	�  J�  	"�  Rn  	t�  S�   	�w  T�   	؜  Y�   	q�  [�  	Ƚ  ^n  	�  _�   	�y  `�   	b�  c�   	+�  f�  	��  i�  	֘ l�   	�J  x�   	��  y�   	ks  �   	�  ��   	J�  ��   	�i  ��   	��  ��  	��  ��  	��  ��  	<� ��  	��  ��  	��  ��  	5�  ��  	<m  ��   	 K  ��   	�R  ��   	op  ��   	�m  ��   	D  ��   	X�  ��   	If  ��   	� ��   	��  ��  	�U  ��  	`  ��  	J�  ��  	��  ��  	� ��  �.  �2  =    	�  �z2  �  �2  =    	� ��2  "  �2  =   	 	,�  ��2  	R�  ��2  "  "  �2  =    	�u  ��2  	��  �0  	�e  ��   �   %3  =   � 	(�  �3  	�  ��   ��  �   �v  �    n�  �    4�  �    *b �    ��  A  	��  ��   	�\  ��  	�  ��3  �  	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  �.  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   (	j4  � *�   �� +�   � ,F4  G /j4  C	�4  x E�   y F�   �{ H�4  (T	�4  `e Vx   x W�  y X�  z Y�    	�  [�4  �a	�5  = c�   F�  d�  �~ eI  h�  fI  
t�  gI  �k hI  tag iI  �N  l
�   ��  o�.  ��  r
�.   iK  u�4  0��  x
�   XS�  {�.  `��  ~R   h��  ��   pu| ��6  x �}  X��6  v1 �A7   v2 �A7  dx ��  dy ��  �  �I  �k �I  tag �I  �W  ��  �o �G7  $��  �57  4SX  ��6  8d�  ��6  @��  �
�   H��  �R   P �6  �5  �z ��4  �	�6  2�  ��   ]  ��  �h  �I  �N  �I  
�K  �I  >} ��6   �6  �}  ��6  
K   �57  ��   �  o�  ��   ��  �7  �4  �  W7  =    �u  ��5  �z �@,  8�	�7  v1 �A7   v2 �A7  82  ��  Mp �y  [�  ��7   �  ��7   SX  ��6  (d�  ��6  0 7  W7  A{ �o7  4	P8  %x �   %y 	�  %dx 
�  %dy �  �o P8  )�  �  0 �  f8  =   =    (} �7  �  *�  &v  @259  @�  459   %x1 5�   %x2 6�   .]  8�  5]  9�  �� :�  ��  =�   �  @�   ��  C�  $�n  G;9  (9x  H;9  0�^  I;9  8 �7  I  >�  K�8  &�h  PR*:  s�  U*:   �H  V*:  %x1 X�   %x2 Y�   %gx \�  %gy ]�  %gz `�   %gzt a�  $�x  d�  (� f�  ,~�  i�  0t  k�  4.� l�   8�  p0:  @	�  r�   H N9  s8  �h  tN9  �	x:  �c  ��   �O  �x:  �x  �
�:   I  �:  =    �  �:  =    I�  �C:  �	�:  �  ��    �  ��:   �:  �  ��:  '��	�;    ��   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  %top �	�;  (��  �	�  U(��  �	�  V(� �	�;  W(�  �	�  � �  �;  =   ? ��  ��:  	.L  &�;  �  	׮  )�;  	�  +�;  	�  ,�;  	�Q  .0:  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7%<  �   	��  8%<  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u Fs<  �:  	��  H�   	��  IA7  	��  K�   	a� L59  	w�  N�   	P{ O�6  	��  Q�   	��  R�<  c7  	��  T�   	�� U�<  f8  	�}  W�   	u| X�7  	M�  Z�   	P�  [�7  	��  a�  	��  b�  	�  c�  	�p  ey  	�T  fi=  �.  	�a  jy  �   �=  =   � 	ը  l{=  y  �=  =   @ 	�p  m�=  	 �  p�  	p|  qy  	$Y  v�   	�K  y�   	g  {�=  �;  	d�  |�=  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   0:  �>  =   =   / 	��  E�>  0:  �>  =   / 	Ԁ  F�>  0:  �>  =   =    	7� G�>  	�R  I�   	��  J0:  	��  U�   	P�  \5  	��  ]5  	L�  ^5  	ߵ  _5  	�  a5  	@�  59  	[�  �7  	 �  �7  	SX  �6  	d�  �6  	��  �   	_�   �   	��  "�  	��  %�  	'�  &�  	�]  (�  A9  �?  =   � 	�P  *�?  	ӯ  +�?  A9  	|  -@  0:  	��  .@  	��  /@  5@  E@  �   �    	��  ;9  �   /@  	qY  "Q@  	�  #Q@  I  �@  =   ? 	��  %u@  	��  &u@  �  �@  =   � 	@Y  (�@  �  �@  =   ? 	V�  )�@  6:  �@  =    	�h  �@  	�  �@  6:  	�  6:  	�f  !u@  	r�  "u@  	��  %;9  	��  &;9  	׆  '�  	��  (�  	�  *�  	��  +�  	�  0:  	��  �   	�_  �   	�_  �   	b  �  	t  �  	j�  ".  	�  :�   	��  ;�   	��  <�   	�W  >0:  	hn  @�  	U~  A�  	�  B�  	 �  C�  	%�  F.  	�u  H.  	z  I.  	- �   	_   �   )�?  '
	��i     )�?  *
	`�i     )�?  +
	��i     *�� -
�  	X�i     *�h  .�   	h�i     *�N  /�   	\�i     *�K  0�   	|�i     )�=  3
	 �i     )�=  5	(�i     )�?  :	H�i     )�?  ;	�i     *D� <
y  	�i     *͊ =
�  	l�i     )�=  >
	d�i     *� ?
�  	��i     *�� @
�  	8�i     *�� A
�  	p�i     *� B
�  	t�i     *щ C
�  	x�i     *S� E�   	D�i     *� F�   	�i     *&� G�   	@�i     *�� H�   	�i     *׊ J
�  	��i     *ߊ K
�  	<�i     *� L
�  	�i     *�� M
�  	L�i     *�� O
�  	$�i     *� P
�  	T�i     *Ɖ R
�  	 �i     *9� S
�  	P�i     *� V@  	�i     *�^  X	;9  	0�i     +_� t��A     {      ��F  ,' u�   T� L� ,�� v�   �� �� -hyp x�  `� \� .|� y�  /� zy  �� �� /� zy  �� �� .\� {�  /0� |�   � � 0�A     �H  �E  1U	?�B     1Ts 1Q|  2K�A     �H  0e�A     �H  !F  1U��� 2��A     �H  2ԮA     �H  0{�A     �H  VF  1U��� 2��A     �H  2��A     �H  2ȳA     �H  2�A     �H  24�A     �H  2S�A     �H  2{�A     �H  2��A     �H  2ƴA     �H  2�A     �H  2��A     �F   3�� ���A           ��G  4Mp �y  5�8 �K   .� (� 6yl ��   �� �� 6yh ��   �� �� 6mid ��   � � 5� ��  H� F� 6top ��   o� k� 5� ��   �� �� 2��A     �H  0��A     I  �G  1T}  0��A     I  �G  1T}  7%�A     I  1T}   8�� `��A           ��H  9ds a�?  �� �� 9x1 b�   M� I� 9x2 c�   �� �� 5�8 eK   �� �� 6col f�H  _� [� 50� g
�   �� �� 5�� h
�   �� �� 2.�A     �H  0b�A     I  �H  1Us  2k�A     I   v4  :��  ��  7:� � :d  d  "	:�� �� �	:�� �� E:�� ��  :�� �� . B6   �  S#  � �*  +�A            �o ��  t�   B   1   int �)  �U   ,	  ^&  �  �1  @�   Q  �    �   	I   62  #	I     &	I   �5  )	I    �@  ,	I   (.  -	I   0*  2B   8;:  5B   < 	�   1  �K 8"l   
�  K  	�   
�  L  
�  M  0t  >  e2    �0  }  ��  2  c   J�  D   �C  
D  ���� �C  Nf  ڵ  RZ  �  c   Y�  ��   �c  |  ��  l  ��  �   c   k1  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {�  c   �p  &�   �  º  GY  �f  ��   v�  �=  c   ��  GQ   ϼ  �  �_  X  &�  �b   �p  	#�  	�  �   S�  	$�  	�  �  j    T}  	%�  	�    j   j    	'	;  acv 	)�  ��  	*�  ��  	+�   �y 	-  �Y  	6;  ��  	:�  s�  	<�   �H  	=�  xz  	>G   	S  x 	@S  =   �  U   �' �  
��  
1�  
]  
4�  	=   =   �  U   � �  
Zy  
8�  �    U   U   � �  
��  
;  Ʃ  
Qc     #  9  U     (  
�  
W9  S  Z  U    E  j  U    
�	�  x �S   y �S  Mp �S  *� �S  ޽  �S   ~x �j  c     @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  c   ��!  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u  (x	"  �u z   � {	B   s |	B   � ~;  N�  �!  ��  �	B   ��  �	B     J]  ��!  "  9"  U   � �^  �("  �   Q"   �  �F"   c   ��%  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  ^"  \	'  �Y  	B    *O  	B   ��  	B   �  	B   b�  	B   ��  	B   �  	B   +�  	B   Zp  	B    o�   	B   $m�  !	B   (4�  "	B   ,�  #	B   0�  $	B   4��  %	B   8L� &	B   <��  '	B   @  (	B   D��  )	B   H\q *	B   Lz�  +	B   P�  ,	B   T/�  -	B   X ʤ  /�%  '  !'  U   � ��  1'  �]  ��)  `e ��   x �1   y �1   z �1    ��  �)  (cN  �)  0Mp �  8�u �  <� �B   @�H  �)  Hr�  �)  P��  �?)  X��  �1   `m�  �1   d��  �1   h  �1   l3F  �1   p8F  �1   t=F  �1   x��  �B   |*� ��%  �y� �E)  �s �B   ��� �K)  ��  �B   ��  �B   �ʺ  �B   ��l  �B   � �  )  ���  B   ���  	B   ��R  ++  �f�  B   �I}  �  ���  )  � 	.'  Gx  �?)  >} ��.   �}  �S  �|  �S  
 	
)  	'  	"  !d  HN++  mo PI-   ��  Q%3  cmd R�2  �  W1   (_  Y1    #_  [1   $bob ]1   (�  aB   ,�[  bB   0sb  dB   4d]  g13  8�W  hA3  P��  i�  h�� lO-  l�N  m1  |E�  p1  ��W  rQ3  �~�  sO-  �*� tO-  ��� wB   ���  xB   �X�  |B   ��e  B   ���  �B   �g  �B   ��u  �B   �|G ��   �Q  �B   ��  �B   �o�  �I-  �"�R  �B    "��  �B   "�  �B   "h  �a3  "I�  ��  @ 	Q)  �z .'  	�  
��  ��   
�\  ��  
�  �h+  �  
��  �B   
��  �B   
2�  ��  
��  �B   
Ɇ  �>+  
��  �B   
��  �B   
�h  �B   
rK  �B   
l�  �B   
]�  �B   
��  �B   C	,  x E1    y F1    �{ H�+  (T	c,  `e V�   x W1   y X1   z Y1     	�  [+,  �a	I-  = c1    F�  d1   �~ eS  h�  fS  
t�  gS  �k hS  tag iS  �N  l
B   ��  oI-  ��  r
O-   iK  uc,  0��  x
B   XS�  {I-  `��  ~j   h��  �B   pu| �.  x 	1+  B   _-  U    �}  X�.  v1 ��.   v2 ��.  dx �1   dy �1   �  �S  �k �S  tag �S  �W  �J  �o ��.  $��  ��.  4SX  ��.  8d�  ��.  @��  �
B   H��  �j   P 	%.  	_-  �z �o,  �	�.  2�  �1    ]  �1   �h  �S  �N  �S  
�K  �S  >} ��.   	+.  �}  �7.  c   ��.  ��   �  o�  ��   ��  ��.  	,  1   �.  U    �u  �_-  �z �
)  8�	r/  v1 ��.   v2 ��.  82  �1   Mp �  [�  �r/   �  �x/   SX  ��.  (d�  ��.  0 	�.  	�.  A{ �/  4	�/  #x 1    #y 	1   #dx 
1   #dy 1   �o �/  )�  Z  0 1   �/  U   U    (} �/  �  *�  	~/  	0  �	T0  �c  ��   �O  �T0  �x  �
d0   S  d0  U    �  t0  U    I�  �0  �	�0  �  �B    �  ��0   	t0  �  ��0  $��	e1    �1    �  �	B   t�  �	B   ��  �	B   /�  �	B   �  �	�  #top �	e1  %��  �	�  U%��  �	�  V%� �	e1  W%�  �	�  � �  v1  U   ? ��  ��0  	�1  ~�  p   �S  
B   ��   
B     !
B   �g  "
B   �^  #
B    ��  %�1  �1  �1  U    
S�  '�1  c   7$2  {�   U�  ~�   >	`2  �� @K)   s A
B   sx B1   sy C1    Nz E$2   	�2  ��  "L   E�  #L  e% $S  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	B   a  2
�  �T  3
�   Mx 4l2  c   1%3  ��   ��  ��   �y  93  B   A3  U    �  Q3  U    �  a3  U    `2  q3  U    hy �Q)  
.L  &�3  	1   
׮  )�3  
�  +�3  
�  ,�3  
�Q  .0  
��  0B   
��  1B   
(_  2B   
դ  4B   
�j  7�3  	B   
��  8�3  
@�  <B   
�O  =B   
(g  >B   
�^  EB   
�u FI4  	�0  
��  HB   
��  I�.  
��  KB   
a� L0  
w�  NB   
P{ O�.  
��  QB   
��  R�4  	�.  
��  TB   
�� U�4  	�/  
�}  WB   
u| Xx/  
M�  ZB   
P�  [r/  
��  a1   
��  b1   
�  c1   
�p  e  
�T  f?5  	q3  
�a  j  B   b5  U   � 
ը  lQ5    5  U   @ 
�p  mn5  
 �  p1   
p|  q  
$Y  vB   
�K  yB   
g  {�5  	v1  
d�  |�5  
- B   
_   B   &4�  %B   	��i     '�5  &	��i     '�5  '	��i     ('� /+�A            � �S   @�  S#  �� �*  6�A     �      �s ��  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  9�  0t  4  e2    �0  }  ��  (  
K   J�  D   �C  
D  ���� �C  N\  ڵ  RP  �  	"|  *�  	��  +�  	I�  ,�  	�a  -�  
K     7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
K   /Q  ��   [r  �4 #�  �   �X  5$  
K   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K]  
�   P�  =_  ��   R�  N�  ��  ��   �p  W�  
K   	32  ��   ({  ��  ğ   F]  	8  
K   	Yw  ��   �c  |  ��  l  ��  �   
K   	k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  	{w  
K   	�  &�   �  º  GY  �f  ��   v�  	��  
K   	�L  GQ   ϼ  �  �_  X  &�  �b   
 	�  ��  
"B   E�  
#B  e% 
$I  u  
%
�  �8 
&
�  ��  
)
�  /b  
-
�  ��  
.	�   a  
2
�  �T  
3
�   Mx 
4L  �  
K   "0  ��  WH  �~  �O  �m  ��   �  ��  ��  	 =� <  ��  .q  ^�  2�   }�  7  �� ;K    	�  r�  �   .� $�  O� )�   �  �  �    0  �  �  �   �  1   �  �  K   R   1    �  ��  ,q  �  �  oS  '  dS  ()r  � +
r   � ,�  @�  -
�   >z .
�   �  /R   �H  3�    �   �  =    
  	�� 7�  	�� 8K   t�   �   �  �  �  =   �' �  	��  1�  	]  4�  �  �  �  =   � �  	Zy  8�  �    =   =   �   	��  ;  Ʃ  QK   .  :  P  =     ?  	�  WP  �p  #m  s  z   S�  $�  �  �  R    T}  %�  �  �  R   R    '	�  acv )a  ��  *z  ��  +�   �y -�  �Y  6�  ��  :4  s�  <4   �H  =4  xz  >�   �  x @�  I  V  =    ;  f  =    
�	�  x �I   y �I  Mp �I  *� �I  ޽  �I   ~x �f  
K   
  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  
K   ��%  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u  (x	&   �u z
    � {	�    s |	�    � ~�   N�  �%   ��  �	�    ��  �	�     J]  ��%  &  5&  =   � !�^  �$&  �   M&  " !�  �B&  #K   ��)  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  Z&  \	 +   �Y  	�     *O  	�    ��  	�    �  	�    b�  	�    ��  	�    �  	�    +�  	�    Zp  	�     o�   	�   $ m�  !	�   ( 4�  "	�   , �  #	�   0 �  $	�   4 ��  %	�   8 L� &	�   < ��  '	�   @   (	�   D ��  )	�   H \q *	�   L z�  +	�   P �  ,	�   T /�  -	�   X ʤ  /�)   +  +  =   � !��  1+  
K   p
,  �! 9& +! v( %# 0  B& @�! ��"  w#  	$  �-  S%  �)   0  @&  ��"    !0    m0    b-    �.    �$     /   @ %   � <"    U-    5'    	!  �]  ���-  `e �:   x ��  y ��  z ��   ��  ��-  (cN  ��-  0Mp �.  8�u �
  <� ��   @�H  ��-  Hr�  ��-  P��  �.  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� ��)  �y� �!.  �s ��   ��� �'.  ��  ��   ��  ��   �ʺ  ��   ��l  ��   �  �  �-  � ��  �   � ��  	�   � �R  0  � f�  �   � I}  �  � ��  �-  � 
,  Gx  �.  >} �4   �}  �I  �|  �I  
 �-   +  &  $d  HN0  mo P�2   ��  Q�9  cmd R�  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g�9  8�W  h�9  P��  i�  h�� l�2  l�N  m�  |E�  p�  ��W  r�9  �~�  s�2  �*� t�2  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��2  �%�R  ��    %��  ��   %�  ��   %h  ��9  %I�  ��  @ -.  �z 
,  	��  ��   	�\  ��  	�  �>0  �  	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  �  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   (	 1  ��  I      I  Vd  !I  �  "I  �� # 1   �   01  =    � %�0  (	`1  � *�   �� +�   � ,<1  G /`1  C	�1  x E�   y F�   �{ Hx1  (T	�1  `e V:   x W�  y X�  z Y�    	�  [�1  �a	�2  = c�   F�  d�  �~ eI  h�  fI  
t�  gI  �k hI  tag iI  �N  l
�   ��  o�2  ��  r
�2   iK  u�1  0��  x
�   XS�  {�2  `��  ~R   h��  ��   pu| ��3  x 0  �   �2  =    �}  X��3  v1 �M4   v2 �M4  dx ��  dy ��  �  �I  �k �I  tag �I  �W  �F  �o �S4  $��  �A4  4SX  �4  8d�  �4  @��  �
�   H��  �R   P �3  �2  �z ��1  �	4  2�  ��   ]  ��  �h  �I  �N  �I  
�K  �I  >} �4   �3  �}  ��3  
K   �A4  ��   �  o�  ��   ��  �4  �1  �  c4  =    �u  ��2  �z ��-  8�	�4  v1 �M4   v2 �M4  82  ��  Mp �.  [�  ��4   �  ��4   SX  �4  (d�  �4  0 4  c4  A{ �{4  4	\5  &x �   &y 	�  &dx 
�  &dy �   �o \5   )�  V  0 �  r5  =   =    (} 5  �  *�  'v  @2A6   @�  4A6   &x1 5�   &x2 6�    .]  8�   5]  9�   �� :�   ��  =�    �  @�    ��  C�  $ �n  GG6  ( 9x  HG6  0 �^  IG6  8 �4  I  >�  K�5  '�h  PR67   s�  U67    �H  V67  &x1 X�   &x2 Y�   &gx \�  &gy ]�  &gz `�   &gzt a�  $ �x  d�  ( � f�  , ~�  i�  0 t  k�  4 .� l�   8 �  p<7  @ 	�  r�   H Z6  5  �h  tZ6  �	�7   �c  ��    �O  ��7   �x  �
�7   I  �7  =    �  �7  =    I�  �O7  �	�7   �  ��     �  ��7   �7  �  ��7  (��	�8     ��    �  �	�    t�  �	�    ��  �	�    /�  �	�    �  �	�  &top �	�8  )��  �	�  U)��  �	�  V)� �	�8  W)�  �	�  � �  �8  =   ? ��  ��7  	9  ~�     �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�8  9  '9  =    	S�  '9  
K   7T9  {�   U�  ~�   >	�9  �� @'.   s A
�   sx B�  sy C�   Nz ET9  
K   1�9  ��   ��  ��   �y  9�9  �   �9  =    �  �9  =    �  �9  =    �9  	:  =    hy �-.  (�	y:  in ��   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�2  �a  �
�   $ ��  �:  ��	;  2�  �
�    I�  ��  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  �;  ( y:  .;  =    ޴  ��:  	.L  &F;  �  	׮  )F;  	�  +F;  	�  ,F;  	�Q  .<7  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�;  �   	��  8�;  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F<  �7  	��  H�   	��  IM4  	��  K�   	a� LA6  	w�  N�   	P{ O4  	��  Q�   	��  Rl<  o4  	��  T�   	�� U�<  r5  	�}  W�   	u| X�4  	M�  Z�   	P�  [�4  	��  a�  	��  b�  	�  c�  	�p  e.  	�T  f�<  	:  	�a  j.  �   =  =   � 	ը  l=  .  <=  =   @ 	�p  m+=  	 �  p�  	p|  q.  	$Y  v�   	�K  y�   	g  {�=  �8  	d�  |�=  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   <7  <>  =   =   / 	��  E&>  <7  X>  =   / 	Ԁ  FH>  <7  z>  =   =    	7� Gd>  	�R  I�   	��  J<7  	��  U�   	P�  \�  	��  ]�  	L�  ^�  	ߵ  _�  	�  a�  	@�  A6  	[�  �4  	 �  �4  	SX  4  	d�  4  	��  �   	_�   �   	��  "�  	��  %�  	'�  &�  	�]  (�  M6  z?  =   � 	�P  *j?  	ӯ  +�?  M6  	|  -�?  <7  	��  .�?  	��  /�?  �?  �?  �   �    	��  G6  �   �?  	qY  "�?  	�  #�?  I  @  =   ? 	��  %@  	��  &@  �  A@  =   � 	@Y  (1@  �  ^@  =   ? 	V�  )M@  B7  z@  =    	�h  j@  	�  �@  B7  	�  B7  	�f  !@  	r�  "@  	��  %G6  	��  &G6  	׆  '�  	��  (�  	�  *�  	��  +�  	�  <7  	��  �   	�_  �   	�_  �   	b  �  	t  �  	j�  "  	�  :�   	��  ;�   	��  <�   	�W  ><7  	hn  @�  	U~  A�  	�  B�  	 �  C�  	%�  F  	�u  H  	z  I  �  	��   M�  	(h   N�   	l�   N�   	�  !.�  	�  !/�  	�  !0�  	�  !2�  	w�  !8Q  	�  !9  	�  !:�  	�_  !;�   	��  !>�  	�  !J�  	"�  !R�  	t�  !S�   	�w  !T�   	؜  !Y�   	q�  ![�  	Ƚ  !^�  	�  !_�   	�y  !`�   	b�  !c�   	+�  !f�  	��  !i�  	֘ !l�   	�J  !x�   	��  !y�   	ks  !�   	�  !��   	J�  !��   	�i  !��   	��  !��  	��  !��  	��  !��  	<� !��  	��  !��  	��  !��  	5�  !��  	<m  !��   	 K  !��   	�R  !��   	op  !��   	�m  !��   	D  !��   	X�  !��   	If  !��   	� !��   	��  !��  	�U  !��  	`  !��  	J�  !��  	��  !��  	� !�2  	:  nD  =    	�  !�^D  �  �D  =    	� !�zD  �  �D  =   	 	,�  !��D  	R�  !��D  �  �  �D  =    	�u  !��D  	��  !�.;  	�e  !��   �   	E  =   � 	(�  !��D  	�  !��  !��  !2  !�v  !�   !n�  !�   !4�  !�   !*b !�   !��  !�A  *�@  D
	�i     *�@  E
	��i     +ϋ G�?  	��i     *�@  K	@�i     *�@  L	��i     *�;  U	x�i     *�;  V	��i     �7  F  =    +s� X�E  	�i     +�� Y�   	ȴi     +A� Z�   	��i     ,z@  	��i     ,�@  	�i     -� �   	شi     -v� >B7  	��i     ,�@  Q		p�i     ,�@  R		дi     ,�@  T
	��i     ,�@  U
	�i     ,�@  	 �i     .�� C@  	@f     .n� D@  	��e     />� ���A     q       ��G  0spr ��@  �� �� 0ds ��?  � � 1��A     �H  2��A     �G  �G  3Us  2��A     �S  �G  3Us  4��A     WI   /� Eu�A           ��H  5spr E!�@  ]� U� 0ds G�?  �� �� 0x H�   �� �� 0r1 I�   %� #� 0r2 J�   J� H� 6� K�  q� m� 6{� L�  �� �� 6��  M�   �� �� 2+�A     �S  �H  3Uv 3Ts 3Q}  1G�A     �S  7��A     vN  3U�U  /� ��A     �       �WI  0i �   z� t� 6r� �   �� �� 0ds �@  	� �� 6< �@  }� {� .�� B7  ��6� �  �� ��  /.� ���A     �       ��I  0i �
�   �� �� 60� �
�   2� 0� 0psp ��I  a� U� 2r�A     �I  �I  3Us� 4��A     �I   �9  /�� ~�A     �      �BK  5psp ~�I  �� �� 0tx ��  C� A� 0x1 ��   h� f� 0x2 ��   �� �� 6� �<  �� �� 6� ��7  �� �� 6�O  ��   ?� =� 6�x  ��  l� j� 0vis ��@  �� �� .K� �B7  ��~29�A     �S  �J  3U	��B      2g�A     �S  K  3U	�B      2��A     �S   K  3Us  1ۿA     �S  8��A     vN  3Uw   /O� ]��A     j       ��K  5sec ]4  �� �� 6�p _�2  � � 60� `�   2� 0� 8�A     �K  3Us   /L� ��A     �      �vN  9�p ��2  [� U� 6�� ��  �� �� 6!� ��  �� �� 0gxt ��  �� �� 0gyt ��  _� [� 0tx ��  �� �� 0tz ��  �� �� 6� ��  �� �� 0x1 ��   3� 1� 0x2 ��   Z� V� 6� �<  �� �� 6� ��7  �� �� 6�O  ��   �� �� 0rot �K   � � 6�x  ��  ?� ;� 6�8 ��   {� w� 0vis ��@  �� �� 0ang �.   � �� 6e  ��  )� #� 25�A     �S  wM  3Us  2F�A     �S  �M  3U}  1h�A     �S  2w�A     �S  �M  3Us  2��A     �S  �M  3U}  2��A     �S  �M  3U	��B      2�A     �S  
N  3U	�B      1�A     �S  2L�A     �S  5N  3Us 3Tv  2z�A     �S  MN  3Tv  1��A     �O  8�A     �S  3U@<$3Tv   /�� ��A     !      �wO  5vis ��@  {� u� 5x1 �	�   �� �� 5x2 �	�   � � 6� �wO  E� A� 6� ��   �� �� 6{q ��  � � 6.� �}O  F� B� 2��A     �S  =O  3T8 1��A     �S  2ѻA     �S  iO  3U	��B      1�A     �O   l1  01  :�� W�A     �       ��O  9� W$wO  �� |� 6×  Y
�   �� �� 6܋ Z
�   +� #� 6P� [�  �� ��  ;2� @�@  ��A     !       �<�� 5�A            �/0{ #ҹA            ��P  9�� #�P  �  � 0i %
�   C� =� 4�A     �P   �   =�� �x�A     Z      �GR  >�� ��P  �� �� ?Wy ��P  �� �� @i �
�   8� 0� @l �
�   �� �� ?� �
�   �� �� ?B� �
�   Z� N� ?' �
�   �� �� @end �
�   /� +� ?ǋ �
�   p� n� 2��A     �S  wQ  3T13Qs  2H�A     �S  �Q  3U~ 3Q4 2x�A     �S  �Q  3U~  2��A     GR  �Q  3R0 2��A     GR  �Q  3U| 3R1 22�A     �S  R  3U	K�B     3Q}�  2e�A     �S  .R  3U	{�B     3Q��� 8��A     �S  3T13Q0  =_� d6�A     B      ��S  >�O  e�   �� �� >� fK   � � >B� gK   j� d� >&� h�  �� �� @r j
�   � � 2f�A     �S  �R  3U	_�B     3T|  2��A     �S  S  3U	��B     3Qv�  2��A     �S  8S  3U	��B     3Qv�  2�A     �S  ^S  3U	��B     3Qv�  8I�A     �S  3U	�B     3Qv� 3R~0  A�� �� "Aɇ ɇ mA��  ��  #7Ad  d  "	AH_  H_  #	Aw� w� sA� � BA� � 6A� � $A�{ �{ = �   �  S#  �� �*  ��A     l      #� x�  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"R   �  K  �   �  L  �  M  9�  0t  2  e2    �J K   �0  }  ��  &  K @  ڵ  RZ  q� �  �� \�  	h0 f   	h1 f  	h2 f  	h3 f  	h4 f  }	 f  	buf 
�  r� 	�   X 
r    =   ? �� ;A�A            �q  �� ;(q  I� C� str ;7�   �� �� ]�A     �  U�UT�T  ~  M� /#�A            ��  �� /'q  �� �� val /=K   �� �� buf 1
�  �l<�A     �  U�UT�lQ4  
r    =    -� �*�A     �       ��  j� ��  :� 4� hd �7q  �� �� t �f  �� �� msb �f  t� r� lsb �f  �� �� p ��  3� � C�A     �  �  Us T0Q0 ��A     �  �  Us T0Q0 ��A     �  Us Tv   r  ^� �H�A     �       ��  hd �"q  -� '� �� �,�  �� y� �� �:1   \� J� j�A     �  n  Us Ts ��A     �  �  Us T0Q0 ��A     �  Us T~ } @  �� 7��A     +      ��  hd 7'q  *  &  "8 71�  n  b  a 9f  D �  b 9f  � G c 9f  � o d 9f  � h e 9f  O � tm 9f   � x :�  ��*�A     )       i G�   <5 :5 p2 H�  h5 `5   
f  �  =    � (�A     ,       �hd ( q  U  �   ��  S#  �� �*  � Q�  ,	  int ^&  9�  e2    �  �0  }  ) n   J @�   � "�    � '
  �� *	(   
 -  �9 0	(    Ml  3	(   $	
 8	(   (C� ;	(   ,� ?	(   0� B/   8   1  	    
!    b    H	_  � K�    C� N	(   "8 Q/   t T/    . V!  : �(   3 �(   � �(   � �(   O �(   �
 ��   	b   �   R �  	_  �   � �  M   r�  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m �  "	�~e     �  t	@ce      L%   ��  S#  �� �*  ]�A     E       Y� p�  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int 	�   �K 8"T   
�  K  �   
�  L  
�  M  9�  0t  9  e2    �0  }  ��  -  K   J�  D   �C  
D  ���� �C  Na  ڵ  RU  	�  K   ��  &�   �  º  GY  �f  ��   v�  ��  	9  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�  9  U  =    
S�  'E  t�  	 �   	a  m  �  =   �' 	r  
��  
1�  
]  
4�  m  m  �  =   � 	�  
Zy  
8�  �  �  =   =   � 	�  
��  
;�  Ʃ  
QK   	�  �    =     	   
�  
W  �p  #.  4  ;   S�  $G  M  X  R    T}  %d  j  z  R   R    '	�  acv )"  ��  *;  ��  +X   �y -z  K     @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  K   ��   �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u  (x	!  �u z   � {	�   s |	�   � ~�  N�  �   ��  �	�   ��  �	�     J]  ��   !  0!  =   � �^  �!  �   H!   �  �=!  \	�"  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /U!  �"  �"  =   � ��  1�"  �   �"  =    (�	@#  in ��   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�"  �a  �
�   $ ��  ��"  ��	�#  2�  �
�    I�  ��  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��#  ( @#  �#  =    ޴  �L#  
�  �   
q  $  �   �   /$  =    	$   �� !/$  $   K   x   Z   �   �   �      �    Ԑ '/$  $   Z   x   x   Z   �   x   x     �#  �$  =    !�� 9�$  	�f     !�� :�   	�f     "ː W��A            �#m- M]�A     D       �=%  $�� M =%  �5 �5 %k�A     C%  &U	�ZB       �#  '?J ?J +	 �G   ��  S#  D� �*  ��A     �      q� ��  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �  	"|  *y  	��  +y  	I�  ,y  	�a  -y  
K   Y�  ��   �c  |  ��  l  ��  �   
K   kP  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {�  
K   ��  &�   �  º  GY  �f  ��   v�  �\  
K   ��  GQ   ϼ  �  �_  X  &�  �b   
K   	"  ��  WH  �~  �O  �m  ��   �  ��  ��  	 (
	d  ��  
B     
 B  Vd  
!B  �  
"B  �� 
#d   �   t  =    � 
%  �   �  =    	N�  %�  	��  '�  �  t   	@  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�  R  =� _  ��  .�  ^�  2!   }�  7�  �� ;K    	�  r�  �   .� $�  O� )   �  �  �    S  �  �  �   �  1     �  K   R   1    �  ��  ,�    oS  '3  dS  ()�  � +
�   � ,�  @�  -
�   >z .
�   �  /R   �H  3�    �   �  =    '  	�� 7�  	�� 8K   H#	  � '
   �^  (1    .�  )	�   (o�  -1   0i�  .	�   8��  /
%  < �   %  =    �   5  =    �  0�  	p�  L�  	t�  M5  	K�  N5  	x�  O5  	��  P5  	��  Q5  	r�  R5  5  �  =    	�  S�  	�u  T5  		�  U5  	h�  V5  t�   �   �  �p  #�  �  �   S�  $      R    T}  %(  .  >  R   R    '	l  acv )�  ��  *�  ��  +   �y ->  �Y  6l  ��  :�  s�  <�   �H  =�  xz  >x   �  x @�  �  �  =   �' �  	��  1�  	]  4�  �  �    =   � �  	Zy  8  �  7  =   =   � !  	��  ;7  Ʃ  QK   H  T  j  =     Y  	�  Wj  B  �  =    4  �  =    
�	�  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x ��  
K   ?  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  
K   ��%  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  uK  (x	L&  �u z?   � {	�   s |	�   � ~l  N�  �%  ��  �	�   ��  �	�     J]  ��%  L&  j&  =   �  �^  �Y&  �   �&  !  �  �w&  "K   ��)  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �&  \	5+  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /�)  5+  R+  =   �  ��  1B+  �]  ��5-  `e ��   x ��  y ��  z ��   ��  �5-  (cN  �5-  0Mp �H  8�u �?  <� ��   @�H  �5-  Hr�  �5-  P��  �p-  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� ��)  �y� �v-  �s ��   ��� �|-  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  5-  ���  �   ���  	�   ��R  \/  �f�  �   �I}  �  ���  5-  � _+  Gx  �p-  >} ��2   �}  �B  �|  �B  
 ;-  5+  L&  #d  HN\/  mo Pt1   ��  Q�9  cmd R@  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g�9  8�W  h:  P��  iy  h�� l�  l�N  mP  |E�  pP  ��W  r:  �~�  s�  �*� t�  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �t1  �$�R  ��    $��  ��   $�  ��   $h  �$:  $I�  �y  @ �-  �z _+  	��  ��   	�\  �y  	�  ��/  �  	��  ��   	��  ��   	2�  �y  	��  ��   	Ɇ  ��  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	J0  x E�   y F�   �{ H*0  (T	�0  `e V�   x W�  y X�  z Y�    	�  [V0  �a	t1  = c�   F�  d�  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  ot1  ��  r
�   iK  u�0  0��  x
�   XS�  {t1  `��  ~R   h��  ��   pu| �:2  x b/  �}  X�:2  v1 ��2   v2 ��2  dx ��  dy ��  �  �B  �k �B  tag �B  �W  �{  �o ��2  $��  ��2  4SX  ��2  8d�  ��2  @��  �
�   H��  �R   P @2  z1  �z ��0  �	�2  2�  ��   ]  ��  �h  �B  �N  �B  
�K  �B  >} ��2   F2  �}  �R2  
K   ��2  ��   �  o�  ��   ��  ��2  J0  �  3  =    �u  �z1  �z �;-  8�	�3  v1 ��2   v2 ��2  82  ��  Mp �H  [�  ��3   �  ��3   SX  ��2  (d�  ��2  0 �2  3  A{ �3  4	�3  %x �   %y 	�  %dx 
�  %dy �  �o �3  )�  �  0 �  4  =   =    (} �3  �  *�  &v  @2�4  @�  4�4   %x1 5�   %x2 6�   .]  8�  5]  9�  �� :�  ��  =�   �  @�   ��  C�  $�n  G�4  (9x  H�4  0�^  I�4  8 �3  B  >�  K.4  &�h  PR�5  s�  U�5   �H  V�5  %x1 X�   %x2 Y�   %gx \�  %gy ]�  %gz `�   %gzt a�  $�x  d�  (� f�  ,~�  i�  0t  k�  4.� l�   8�  p�5  @	�  r�   H �4  !4  �h  t�4  �	&6  �c  �y   �O  �&6  �x  �
66   B  66  =    �  F6  =    I�  ��5  �	z6  �  ��    �  �z6   F6  �  �S6  '��	77    ��   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  %top �	77  (��  �	�  U(��  �	�  V(� �	77  W(�  �	�  � �  H7  =   ? ��  ��6  0 	�7  x $
�    y %
�   ��  (	�   �� +
�   num .
�7  on 2�7  p 5�7   "8 8	�   ( �   y  �  �� :U7  8@	�7  n C�7   p F�  0 � H�7  0M	h8  x P�    y Q�   <� T�   ?� W�7  on [�7  p ^�7   "8 a�   ( �� c
8  0j	�8  x m�    y n�   � qy  val t�7  on x�7  p {�   "8 |�   ( � ~t8  	69  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�8  69  R9  =    	S�  'B9  
K   79  {�   U�  ~�   >	�9  �� @|-   s A
�   sx B�  sy C�   Nz E9  
K   1�9  ��   ��  ��   �y  9�9  �   :  =    y  :  =    y  $:  =    �9  4:  =    hy ��-  	.L  &L:  �  	׮  )L:  	�  +L:  	�  ,L:  	�Q  .�5  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�7  	��  8�7  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F;  �6  	��  H�   	��  I�2  	��  K�   	a� L�4  	w�  N�   	P{ O�2  	��  Q�   	��  Rl;  3  	��  T�   	�� U�;  4  	�}  W�   	u| X�3  	M�  Z�   	P�  [�3  	��  a�  	��  b�  	�  c�  	�p  eH  	�T  f�;  4:  	�a  jH  �   <  =   � 	ը  l<  H  <<  =   @ 	�p  m+<  	 �  p�  	p|  qH  	$Y  v�   	�K  y�   	g  {�<  H7  	d�  |�<  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   �5  <=  =   =   / 	��  E&=  �5  X=  =   / 	Ԁ  FH=  �5  z=  =   =    	7� Gd=  	�R  I�   	��  J�5  	��  U�   	P�  \L  	��  ]L  	L�  ^L  	ߵ  _L  	�  aL  	@�  �4  	[�  �3  	 �  �3  	SX  �2  	d�  �2  	��  �   	_�   �   	��  "y  	��  %y  	'�  &y  	�]  (y  �4  z>  =   � 	�P  *j>  	ӯ  +�>  �4  	|  -�>  �5  	��  .�>  	��  /�>  �>  �>  �   �    	��   �4  �    �>  	qY   "�>  	�   #�>  B  ?  =   ? 	��   %?  	��   &?  �  A?  =   � 	@Y   (1?  �  ^?  =   ? 	V�   )M?  �5  z?  =    	�h  !j?  	�  !�?  �5  	�  !�5  	�f  !!?  	r�  !"?  	��  !%�4  	��  !&�4  	׆  !'�  	��  !(�  	�  !*�  	��  !+�  	�  "�5  	��  "�   	�_  "�   	�_  "�   	b  "�  	t  "�  	j�  ""�  	�  ":�   	��  ";�   	��  "<�   	�W  ">�5  	hn  "@�  	U~  "A�  	�  "B�  	 �  "C�  	%�  "F�  	�u  "H�  	z  "I�  	��  (y  )n� 1�  	��i     *�� �y�A     �       ��A  +bi  �A  #6 6 ,"O  y  �6 �6 -x �   �6 �6 -y �   7 7 -w �   +7 )7 -h �   X7 V7 .��A     �G  �A  /U	��B      0��A     �G  1�A     �G  /U|  /Tv�~/R} 0$0&/X~ 0$0&/Y|    �8  *� �`�A            �mB  2b ��A  U2x �	�   T2y �	�   Q2i ��  R2val ��7  X2on ��7  Y *�� ���A     �       �RC  3mi �RC  �7 �7 4"O  �y  �7 �7 5w ��   >8 <8 5h ��   e8 a8 5x ��   �8 �8 5y ��   �8 �8 .�A     �G  C  /U	��B      .0�A     �G  DC  /U| /Tv�~/R} /Y|  0K�A     �G   h8  *[� �{�A            ��C  2i �RC  U2x �	�   T2y �	�   Q2il ��7  R6?� �
�7  X2on ��7  Y * �N�A     -       �3D  3per �3D  �8 �8 4"O  �	�   U9 M9 0q�A     �G  7{�A     $E  /U�U/T�T  �7  *� �+�A     #       �$E  2p �3D  U2x �	�   T2y �	�   Q2pl ��7  R2num �
�7  X2on ��7  Y6� ��  � 8�F  +�A     �  �9G  �9 �9 9�F  �9 �9 9�F  : �9 9�F  &: $: 9�F  K: I: 9�F  p: n: 9�F  �: �:   *�� ��A            ��E  3n ��E  �: �: 4"O  �y  ; 
; 7*�A     �E  /U�U/T�T  �7  *�� T��A     A      ��F  3n U�E  f; \; 4"O  Vy  �; �; :֑ Y
�   5num Z
�   "< < 5w \
�   �< �< 5h ]
�   �< �< 5x ^
�   = = 5neg `
�   ]= Y= .c�A     �G  XF  /U	��B      .��A     �G  vF  /U} /Y}  .��A     �G  �F  /U}   .��A     �G  �F  /U}  ;�A     �G   <M� ;G  =n <�E  =x =	�   =y >	�   =pl ?�7  =num @
�7  =on A�7  >��  B	�    *&� 3��A            �PG  1��A     �G  /U	��B     /T1  ?�F  ��A             ��G  @�F  U@�F  T@�F  Q@�F  R@�F  X@�F  Y@G  �  A��  ��  #7Ay�  y�  9A1� 1� 5A��  ��  C 8m   ��  S#  �� �*  0�A     �      �� I�  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  
K   Jy  D   �C  
D  ���� �C  NU  ڵ  RI  �   	"  ��  ";   E�  #;  e% $B  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4�  
K   ![  �p   �  ��  S�  ��   �F  '.  *	�  *� ,[   "G  C	�   (G  C�   �]  C�   :G  C�    �U  Dg  �  �  	��  	��   	�\  	�y  	�  	��  �  	��  	��   	��  	��   	2�  	�y  	��  	��   	Ɇ  	��  	��  	��   	��  	��   	�h  	��   	rK  	��   	l�  	��   	]�  	��   	��  	��   
K   
"�  ��  WH  �~  �O  �m  ��   �  ��  ��  	 
K     7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
K   /O  ��   [r  �4 #�  �   �X  5"  
K   :�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K[  
�   P�  =_  ��   R�  N�  ��  ��   �p  W�  =�   ��  .J  ^�  2�   }�  7�  �� ;K    	{  r�  �   .� $�  O� )�   �  �  �    	  {  �  �   �  1   �  �  K   R   1    �  ��  ,J  �  oS  '�  dS  ()E  � +
E   � ,�  @�  -
�   >z .
�   �  /R   �H  3U    �   U  =    �  	�� 7U  	�� 8K   	"|  *y  	��  +y  	I�  ,y  	�a  -y  
K   3�  ��   ({  ��  ğ   F]  8�  
K   Y  ��   �c  |  ��  l  ��  �   
K   k`  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {  
K   ��  &�   �  º  GY  �f  ��   v�  �l  
K   ��  GQ   ϼ  �  �_  X  &�  �b   	� M�   	5 N�   H#	T  � '
T   �^  (1    .�  )	�   (o�  -1   0i�  .	�   8��  /
d  < �   d  =    �   t  =    �  0�  
K   :�  ��  u�  � >�  
K   C�  `�  � 0�  Ւ H�  	p�  L�  	t�  Mt  	K�  Nt  	x�  Ot  	��  Pt  	��  Qt  	r�  Rt  t  8	  =    	�  S(	  	�u  Tt  		�  Ut  	h�  Vt  t�   �   h	  �p  #�	  �	  �	   S�  $�	  �	  �	  R    T}  %�	  �	  �	  R   R    '	�	  acv )y	  ��  *�	  ��  +�	   �y -�	  �Y  6�	  ��  :L
  s�  <L
   �H  =L
  xz  >
   
  x @
  t	  o
  =   �' ^
  	��  1o
  	]  4�
  t	  t	  �
  =   � �
  	Zy  8�
  �  �
  =   =   � �
  	��  ;�
  Ʃ  QK   �
  �
  �
  =     �
  	�  W�
  B    =    4  .  =    
�	u  x �B   y �B  Mp �B  *� �B  ޽  �B   ~x �.  
K   �  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��  
K   �e(  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�  (x	�(   �u z�    � {	�    s |	�    � ~�	   N�  e(   ��  �	�    ��  �	�     J]  �r(  �(  �(  =   � !�^  ��(  �   )  " !�  �
)  #K   �n,  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  ")  \	�-   �Y  	�     *O  	�    ��  	�    �  	�    b�  	�    ��  	�    �  	�    +�  	�    Zp  	�     o�   	�   $ m�  !	�   ( 4�  "	�   , �  #	�   0 �  $	�   4 ��  %	�   8 L� &	�   < ��  '	�   @   (	�   D ��  )	�   H \q *	�   L z�  +	�   P �  ,	�   T /�  -	�   X ʤ  /{,  �-  �-  =   � !��  1�-  �]  ���/  `e �R
   x �h	  y �h	  z �h	   ��  ��/  (cN  ��/  0Mp ��
  8�u ��  <� ��   @�H  ��/  Hr�  ��/  P��  �0  X��  �h	  `m�  �h	  d��  �h	  h  �h	  l3F  �h	  p8F  �h	  t=F  �h	  x��  ��   |*� �n,  �y� �	0  �s ��   ��� �0  ��  ��   ��  ��   �ʺ  ��   ��l  ��   �  �  �/  � ��  �   � ��  	�   � �R  �1  � f�  �   � I}  u  � ��  �/  � �-  Gx  �0  >} ��4   �}  �B  �|  �B  
 �/  �-  �(  $d  HN�1  mo P�3   ��  Q=<  cmd R"  �  Wh	  (_  Yh	   #_  [h	  $bob ]h	  (�  a�   ,�[  b�   0sb  d�   4d]  gj<  8�W  hz<  P��  iy  h�� l�3  l�N  m`  |E�  p`  ��W  r�<  �~�  s�3  �*� t�3  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��3  �%�R  ��    %��  ��   %�  ��   %h  ��<  %I�  �y  @ 0  �z �-  (	M2  ��  B      B  Vd  !B  �  "B  �� #M2   �   ]2  =    � %2  C	�2  x Eh	   y Fh	   �{ Hi2  (T	�2  `e VR
   x Wh	  y Xh	  z Yh	    	�  [�2  �a	�3  = ch	   F�  dh	  �~ eB  h�  fB  
t�  gB  �k hB  tag iB  �N  l
�   ��  o�3  ��  r
�3   iK  u�2  0��  x
�   XS�  {�3  `��  ~R   h��  ��   pu| ��4  x �1  �   �3  =    �}  X��4  v1 �>5   v2 �>5  dx �h	  dy �h	  �  �B  �k �B  tag �B  �W  �  �o �D5  $��  �25  4SX  ��4  8d�  ��4  @��  �
�   H��  �R   P �4  �3  �z ��2  �	�4  2�  �h	   ]  �h	  �h  �B  �N  �B  
�K  �B  >} ��4   �4  �}  ��4  
K   �25  ��   �  o�  ��   ��  �5  �2  h	  T5  =    �u  ��3  �z ��/  8�	�5  v1 �>5   v2 �>5  82  �h	  Mp ��
  [�  ��5   �  ��5   SX  ��4  (d�  ��4  0 �4  T5  A{ �l5  4	M6  &x h	   &y 	h	  &dx 
h	  &dy h	   �o M6   )�    0 h	  c6  =   =    (} �5  �  *�  'v  @227   @�  427   &x1 5�   &x2 6�    .]  8h	   5]  9h	   �� :h	   ��  =�    �  @h	    ��  Ch	  $ �n  G87  ( 9x  H87  0 �^  I87  8 �5  B  >�  K}6  '�h  PR'8   s�  U'8    �H  V'8  &x1 X�   &x2 Y�   &gx \h	  &gy ]h	  &gz `h	   &gzt ah	  $ �x  dh	  ( � fh	  , ~�  ih	  0 t  kh	  4 .� l�   8 �  p-8  @ 	�  r�   H K7  p6  �h  tK7  �	u8   �c  �y    �O  �u8   �x  �
�8   B  �8  =    �  �8  =    I�  �@8  �	�8   �  ��     �  ��8   �8  �  ��8  (��	�9     �h	    �  �	�    t�  �	�    ��  �	�    /�  �	�    �  �	�  &top �	�9  )��  �	�  U)��  �	�  V)� �	�9  W)�  �	�  � �  �9  =   ? ��  ��8  0 	:  x $
�    y %
�   ��  (	�   �� +
�   num .
:  on 2:  p 5:   "8 8	�   ( �   y  !:  ]2  �� :�9  8@	S:  n C':   p F!:  0 � H3:  0M	�:  x P�    y Q�   <� T�   ?� W:  on [:  p ^:   "8 a�   ( �� c_:  0j	';  x m�    y n�   � qy  val t:  on x:  p {!:   "8 |�   ( � ~�:  	�;  ~�  �   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %3;  �;  �;  =    	S�  '�;  
K   7�;  {�   U�  ~�   >	<  �� @0   s A
�   sx Bh	  sy Ch	   Nz E�;  
K   1=<  ��   ��  ��   �y  9<  
K   @j<  el �l �l  �   z<  =    y  �<  =    y  �<  =    <  �<  =    hy �0  (�	=  in �y   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�3  �a  �
�   $ ��  ��<  ��	�=  2�  �
�    I�  �y  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��=  ( =  �=  =    ޴  �&=  	.L  &�=  h	  	׮  )�=  	�  +�=  	�  ,�=  	�Q  .-8  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7:  	��  8:  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�>  �8  	��  H�   	��  I>5  	��  K�   	a� L27  	w�  N�   	P{ O�4  	��  Q�   	��  R?  `5  	��  T�   	�� U%?  c6  	�}  W�   	u| X�5  	M�  Z�   	P�  [�5  	��  ah	  	��  bh	  	�  ch	  	�p  e�
  	�T  f�?  �<  	�a  j�
  �   �?  =   � 	ը  l�?  �
  �?  =   @ 	�p  m�?  	 �  ph	  	p|  q�
  	$Y  v�   	�K  y�   	g  {@  �9  	d�  |@  	��    h	  		�   !h	  	�3  #�   	_   $�   	-�   (�   	�f   )�   	�G   +h	  	`�   ,h	  	A�   -h	  	��   /�   	��   1�   	P�   2�   -8  �@  =   =   / 	��   E�@  -8  �@  =   / 	Ԁ   F�@  -8  A  =   =    	7�  G�@  	�R   I�   	��   J-8  	��   U�   	P�   \�  	��   ]�  	L�   ^�  	ߵ   _�  	�   a�  	@�  !27  	[�  !�5  	 �  !�5  	SX  !�4  	d�  !�4  	��  !�   	_�  ! �   	��  !"y  	��  !%y  	'�  !&y  	�]  !(y  >7  B  =   � 	�P  !*B  	ӯ  !+-B  >7  	|  !-?B  -8  	��  !.?B  	��  !/?B  cB  sB  �   �    	��  "87  �  " ]B  	qY  ""B  	�  "#B  B  �B  =   ? 	��  "%�B  	��  "&�B  h	  �B  =   � 	@Y  "(�B  h	  �B  =   ? 	V�  ")�B  38  C  =    	�h  #C  	�  #-C  38  	�  #38  	�f  #!�B  	r�  #"�B  	��  #%87  	��  #&87  	׆  #'h	  	��  #(h	  	�  #*h	  	��  #+h	  	�  $-8  	��  $�   	�_  $�   	�_  $�   	b  $h	  	t  $h	  	j�  $"�  	�  $:�   	��  $;�   	��  $<�   	�W  $>-8  	hn  $@h	  	U~  $Ah	  	�  $Bh	  	 �  $Ch	  	%�  $F�  	�u  $H�  	z  $I�  	ʓ  %CR
  u  �D  =    	��  %b�D  �   �D  =    	��  %c�D  	0K  %d�   	?�  %e�   %�	E  x %�h	   y %�h	  dx %�h	  dy %�h	   ��  %��D  %�9E  �p %�
�3  ��  %�
�5   %�	hE  {q %�h	   ��  %�y  d %�	E   t�  %�9E  hE  �E  =   � 	r %�tE  	�T  %��E  hE  	l�  %�h	  	�  %�h	  	?k  %�h	  	�d  %�h	  	2~ %�E  	��  %�y  	��  %�h	  	k�  %�h	  	Z�  %��5  �5  F  =    	�v  %�F  	�v  %��   	"�  %��3  !�  %�  !�U  %87  !��  %87  !t�  %�   !�  %	�   !.Y  %
h	  !7Y  %h	  !�h  %�F  �3  !*� %�3  !<i  %�3  	G  &y  	��  &�   �   �F  =    
K   &�G  *top  �G  �  �]  &��F   &�	jG  ��  &��5   ��  &�G  O{  &�
�   ��  &�
�   iK  &�jG   �2  ��  &�G  pG  �G  =    	��  &�|G  #K   &�G  *up  �  �F  �S   FT  &
�G  #K   &�G  ��   �x  H�  ��  �H   ��  &�G  H&	�H   `e &R
    >} &�4   L� &h	   &low &h	  $ +� & h	  ( �Z &!
�   , r� &"
�   0 �f  &#�G  4 �f  &$�G  8 ��  &%y  <&tag &&
�   @ *� &'�G  D �w &)H  �H  �H  =    �H  !�  &2�H  #K   &�I  ��   �s  z�  ��  �T  ܭ   gY  &��H  H&�	�I   `e &�R
    *� &�I   >} &��4    �W  &�h	  ( �}  &�h	  , L� &�h	  0 ��  &�y  4 ��  &�
�   8&tag &�
�   < ��  &�
�   @  w &�+I  �I  �I  =    �I  !j�  &�I  	��  '.t  ) (
J  J @(�J  � ("�    � ('
�F  �� (*	�   
 (-�J  �9 (0	�    Ml  (3	�   $	
 (8	�   (C� (;	�   ,� (?	�   0� (BR   8 �I   (H	�J  � (K�    C� (N	�   "8 (QR   t (TR    . (V�J  	: (��   	3 (��   	� (��   	� (��   	O (��   	�
 (��   �I  =K  " 	R )2K  �J  TK  " 	� )IK  
K   )$M  z  � �     & / 8 	; 
D M V _ h q z � q o z � � � � � � _ � o x �  � !�	 "  #1
 $� %< &( 'l
 (: )�	 *� +�
 ,� -V
 .# /� 0V 1� 2� 3� 4� 5a
 6� 7�
 8� 9� :D ;� <� =6 >f ?� @* Aa B C� D 	 *V�   	N�  +%�3  	��  +'�  "  	��  ,My  	(h  ,N�   	l�  ,N�   	�  -.y  	�  -/y  	�  -0y  	�  -2y  	w�  -8O  	�  -9  	�  -:�  	�_  -;�   	��  ->y  	�  -Jy  	"�  -R�  	t�  -S�   	�w  -T�   	؜  -Y�   	q�  -[y  	Ƚ  -^�  	�  -_�   	�y  -`�   	b�  -c�   	+�  -fy  	��  -iy  	֘ -l�   	�J  -x�   	��  -y�   	ks  -�   	�  -��   	J�  -��   	�i  -��   	��  -�y  	��  -�y  	��  -�y  	<� -�y  	��  -�y  	��  -�y  	5�  -�y  	<m  -��   	 K  -��   	�R  -��   	op  -��   	�m  -��   	D  -��   	X�  -��   	If  -��   	� -��   	��  -�y  	�U  -�y  	`  -�y  	J�  -�y  	��  -�y  	� -��  �<  �O  =    	�  -��O  y  �O  =    	� -��O  u  �O  =   	 	,�  -��O  	R�  -�P  u  u  )P  =    	�u  -�P  	��  -��=  	�e  -��   �   ^P  =   � 	(�  -�MP  	�  -�y  !��  -�  !�v  -�   !n�  -�   !4�  -�   !*b -�   !��  -1M  	Y�  .%
)  	��  .&
)  +�  	 �i     ,�  
�?  	`%f     ,�� y  	X%f     ,5� �   	T%f     ,�� K   	P%f     ,�� �   	L%f     -Q� �  -� �  ,�� y  	H%f     -�� "y  ,� %y  	D%f     -H� (y  ,И +y  	@%f     ,�� .y  	<%f     ,�� 1y  	8%f     ,l 4!:  	0%f     !:  0R  =   	 ,�� 7 R  	�$f     ,� :!:  	�$f     ,� = R  	�$f     !:  �R  =    ,�" @uR  	@$f     !:  �R  =   ) ,X� C�R  	�"f     ,� F!:  	�"f     ,�� I!:  	�"f     !:  S  =   =    ,i� L�R  	`"f     ,�� O':  	 "f     ,#� R':  	�!f     ,�� US:  	�!f     ,�� X';  	`!f     �:  �S  =    ,g� \zS  	@ f     ,V� _�:  	  f     �:  �S  =    ,�� b�S  	`f     ,� eS:  	 f     ':  T  =    ,� h�S  	`f     ,(� k�S  	�f     ,2� p�   	�f     ,_� s�   	h�e     ,̜ v�<  	`f     ,L� y�   	Pf     ,:� |�   	Lf     �   �T  =    ,�� �T  	@f     ,Œ ��   	8f     +�  �	 �e     +�  �	��e     +�  �	`�e     +	  �	 �e     +	  �	��e     +	  �	@�e     +8	  �	@�e     +D	  �	��e     +P	  �	��e     +\	  �	 �e     ,~� ��   	4f     � /�U  �U  �U  �   :   ,�� jy  	�e     .J ���A             �@V  /��A     �\  0��A     �k  1U
 (1T11Q0  2� y.t m��A     %       ��V  /��A     @V  /��A     �[  /��A     �V   .�� ���A     �      ��[  3i �	�   �= �= 4&�A     �k  W  1U	 "f     1T,1Q�1R	�$f     1Y	H%f      4a�A     l  MW  1U	�!f     1TZ1Q�1R	�$f     1Y	H%f      4��A     l  �W  1U	`!f     1Th1Q�1X	@%f     1Y	H%f      4��A     l  �W  1U|P1Rs4$`"f     "1Y	<%f      4�A     �k  X  1U	�!f     1T�1Q�1R	�$f     1X	�f     1Y	8%f      4'�A     l  mX  1U	  f     1T�1Q�1R	�"f     1X	Lf     1Y	H%f      4X�A     l  �X  1U	 f     1T�1Q�1R	�$f     1Y	H%f      4}�A     l  Y  1U	`f     1T�1Q�1R	@$f     1X	@f     1Y	H%f      4��A     l  VY  1U	�f     1T�1Q�1R	@$f     1X	Df     1Y	H%f      4��A     l  �Y  1U	�f     1T�1Q�1R	@$f     1X	Hf     1Y	H%f      4��A     �k  �Y  1U	`f     1T
 1Q�1R	�$f     1Y	H%f      4/�A     �k  4Z  1U	�f     1T
 1Q�1R	�$f     1Y	H%f      4c�A     �k  zZ  1U	�f     1T
 1Q�1R	�$f     1Y	H%f      4��A     �k  �Z  1U	�f     1T
 1Q�1R	�$f     1Y	H%f      4��A     �k  [  1U	�f     1T
:1Q�1R	�$f     1Y	H%f      4��A     �k  L[  1U	�f     1T
:1Q�1R	�$f     1Y	H%f      43�A     �k  �[  1U	 f     1T
:1Q�1R	�$f     1Y	H%f      0g�A     �k  1U	0f     1T
:1Q�1R	�$f     1Y	H%f       .l� �F�A     �       �\  3i �
�   �= �= 5��A     'l   .� �D�A            �B\  5F�A     B\   .�� �:�A     
       �}\  6D�A     �]  1U	��A       7�� ���A            ��\  8� �%�   d> `> 8�R �9:  �> �> 0��A     3l  1U�U  .� �&�A            �(]  41�A     ?l  ]  1U	�RB      5:�A     (]   .ח ��A     
       �c]  6&�A     �]  1U	0�A       7�� �0�A            ��]  8� �#�   �> �> 8�R �7:  2? ,? 0>�A     Kl  1U�U1T1  7V� 4C�A     `      �db  8�� 43�U  �? ~? 3i 7
�   �? �? 3j 8
�   �@ �@ 9w� 9
�   6A A ,��  ;
�F  �G4t�A     Wl  v^  1U�G1T91Q	�B     1Rv  :��A     �^  1U�G1T| �$f     " 4��A     Wl  �^  1U�G1T91Q	�B      :��A     �^  1U�G1T| �$f     " :��A     _  1U	%�B     1T	�$f      4��A     Wl  @_  1U�G1T91Q	.�B     1Rv  :��A     f_  1U�G1Tv3$@$f     " :��A     �_  1U	7�B     1T	�"f      4�A     Wl  �_  1U�G1T91Q	>�B     1Rv :.�A     �_  1U�G1T| `"f     " 4k�A     Wl  `  1U�G1T91Q	G�B      :w�A     -`  1U�G1T	�"f      :��A     U`  1U	N�B     1T	0%f      4��A     Wl  �`  1U�G1T91Q	T�B     1Rv 1X} :��A     �`  1U�G1T~x 4��A     Wl  �`  1U�G1T91Q	^�B     1Rv  :��A     �`  1U�G1T| 4��A     Wl  a  1U�G1T91Q	g�B     1Rv  :�A     9a  1U�G1T|  4�A     Wl  ia  1U�G1T91Q	p�B     1Rv  :'�A     �a  1U�G1T|( 4?�A     Wl  �a  1U�G1T91Q	z�B     1Rv  :K�A     �a  1U�G1T|0 4e�A     Wl  �a  1U�G1T91Q	��B     1Rv :u�A     b  1U�G1T|x :��A     ?b  1U	��B     1T	 $f      ;��A     1U	��B     1T	($f       . ��A     A       ��b  8rK  y  �B �B 8"O  -y  �B �B /�A     He  5�A     c  5�A     �b   .�� ��A            �c  6��A     Hc  1U0  .� ��A            �Hc  /��A     k  6��A     Hc  1U1  .o� ���A     �       �He  8"O  �y  �B �B 3i �
�   RC JC 4�A     cl  �c  1U	 "f     1Ts  4�A     cl  �c  1Uv `f     "1Ts  41�A     cl  d  1Uv pf     "1Ts  4K�A     ol  )d  1U	�!f     1Ts  4W�A     ol  Nd  1U	 f     1Ts  4c�A     {l  sd  1U	`!f     1Ts  4q�A     �l  �d  1UvP1Ts  4��A     �l  �d  1U	  f     1Ts  4��A     �l  �d  1U	`f     1Ts  4��A     �l   e  1U	�f     1Ts  4��A     �l  %e  1U	�f     1Ts  6��A     cl  1U	�!f     1T�U  .�� ��A     �       ��e  9@� �
�   �C �C <pal ��  3cnt �
�   9D 3D 3bzc �
�   �D �D 4��A     �l  �e  1T8 5��A     �l   .e$ ���A     )       �f  /��A     �l  /��A     f   .� \��A     �       �if  ,B� ^�   	 �e     3i _
�   
E �D /f�A     if   .L� ��A     �      �qg  3i �
�   �E �E 9R� ��
  �E �E 9�� ��
  
F F ,�� ��   	�e     ,�� ��   	�f     9G� �y  FF @F /��A     qg  /�A     qg  /8�A     �l  /w�A     qg  /��A     qg  /��A     qg  /K�A     qg  /��A     qg   =�� ��   ��A     A       ��g  9�  �
�   �F �F ,2� ��   	�f     ,b� ��   	�e      =Y�  �y  &�A     �      ��j  >ev ��j  �F �F 3i ��   @G G ?��A     �       �h  @buf �j  �]9� �   �H �H 4�A     �l  �h  1U	 �e     1T�] 0~�A     �l  1T1  ?��A     H       �h  @buf Q�j  	 f     0�A     �l  1U	 f     1T41Q	��B       ?&�A     �       ri  @buf ]�j  �]92�  ^�   2I .I 3map _�   mI iI 45�A     �l  di  1U	��e     1T�] /��A     �l   4��A     �l  �i  1U	��e      4��A     �l  �i  1U	��e      4
�A     �l  �i  1U	 �e      4s�A     �l  �i  1U	`�e      4��A     �l  j  1U	 �e      4��A     �l  ,j  1U	@�e      4��A     �l  Kj  1U	��e      4�A     �l  pj  1Uv H@�e     " 4'�A     �l  �j  1Tv  4h�A     �l  �j  1U	��e      4��A     �l  �j  1U	��e      0��A     �l  1U	 �e       �  �   �j  =    �   k  =   3 22� �Ak  ��A     q       ��k  /��A     m  4��A     m  Vk  1U01T0 4��A     m  sk  1U�1T0 /��A     #m  0 �A     /m  1U01T01R
@1X 1Y0  A@V  n�A     /       ��k  4��A     �l  �k  1T8 /��A     �l   B� � 
6BM� M� �B� � �B� � �B[� [� �B&� &� �B�q  �q  J	B�{ �{ =B��  ��  CB[�  [�  fB�� �� �B  �B�� �� �B�� �� �B� � BB� � 	hB� � /BEf Ef  xB,M ,M 9BL L *ABG�  G�  0/B� � &B�~  �~  3B#m #m 1	Bw� w� +RBy�  y�  +9B� � +VB1� 1� +5 [   ;�  S#  r� �*  ��A     �      �� ��  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  9�  0t  4  e2    �0  }  ��  (  
K   J�  D   �C  
D  ���� �C  N\  ڵ  RP  �  ) �  J @9  � "�    � '
9  �� *	�   
 -I  �9 0	�    Ml  3	�   $	
 8	�   (C� ;	�   ,� ?	�   0� BR   8 �   I  =    �   H	�  � K�    C� N	�   "8 QR   t TR    . VO  
K   Y�  �?  N> �> i? �? ~? �? D@ A �? 	�@ 
 �  �  R    �  	: ��   	3 ��   	� ��   	� ��   	O ��   	�
 ��    	�  ��  "B   E�  #B  e% $I  u  %
�  �8 &
�  ��  )
�  /b  -
�  ��  .	�   a  2
�  �T  3
�   Mx 4J  
K   	-  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  	(�  
K   	/f  ��   [r  �4 #�  �   �X  	59  
K   	:�  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  	Kr  
�   	P  =_  ��   R�  N�  ��  ��   �p  	W�  
K   
3G  ��   ({  ��  ğ   F]  
8   
K   
Y�  ��   �c  |  ��  l  ��  �   
K   
k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  
{�  
K   
�  &�   �  º  GY  �f  ��   v�  
��  
K   
�a  GQ   ϼ  �  �_  X  &�  �b   �   q  =    I  �  =    ;  �  =    
�	�  x �I   y �I  Mp �I  *� �I  ޽  �I   ~x ��  �  �   �  �  	��  M�  	(h  N�   	l�  N�   	y  ~�     �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %!  y  �  =    	S�  '�  t�   �   �  �  �  =   �' �  	��  1�  	]  4�  �  �  �  =   � �  	Zy  8�  �    =   =   �   	��  ;  Ʃ  QK   /  ;  Q  =     @  	�  WQ  �p  #�  S�  $�  T}  %�  �  �  R   R    '	�  acv )b  ��  *n  ��  +z   �y -�  �Y  6�  ��  :	  s�  <	   �H  =	  xz  >�   �  x @�  
K   z  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  �)	  
K   �&  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u�  (x	�&  �u zz   � {	�   s |	�   � ~�  N�  &  ��  �	�   ��  �	�     J]  �&  �&  �&  =   �  �^  ��&  �   �&  !  �  ��&  "K   �*  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  �&  \	p+  �Y  	�    *O  	�   ��  	�   �  	�   b�  	�   ��  	�   �  	�   +�  	�   Zp  	�    o�   	�   $m�  !	�   (4�  "	�   ,�  #	�   0�  $	�   4��  %	�   8L� &	�   <��  '	�   @  (	�   D��  )	�   H\q *	�   Lz�  +	�   P�  ,	�   T/�  -	�   X ʤ  /#*  p+  �+  =   �  ��  1}+  
K   7�+  {�   U�  ~�   >	�+  �� @�+   s A
�   sx B�  sy C�   �&  Nz E�+  �]  ���-  `e �	   x ��  y ��  z ��   ��  ��-  (cN  ��-  0Mp �/  8�u �z  <� ��   @�H  ��-  Hr�  ��-  P��  �.  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� �*  �y� � .  �s ��   ��� ��+  ��  ��   ��  ��   �ʺ  ��   ��l  ��   � �  �-  ���  �   ���  	�   ��R   0  �f�  �   �I}  �  ���  �-  � 	,  Gx  �.  >} �=   �}  �I  �|  �I  
 �-  p+  #d  HN 0  mo P@0   ��  Q40  cmd R�  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  gF0  8�W  hV0  P��  i�  h�� lf0  l�N  m�  |E�  p�  ��W  rv0  �~�  sf0  �*� tf0  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  �@0  �$�R  ��    $��  ��   $�  ��   $h  ��0  $I�  ��  @ &.  �z 	,  
K   140  ��   ��  ��   �y  90  0  �   V0  =    �  f0  =    �   v0  =    �  �0  =    �+  �0  =    hy �&.  (�	1  in ��   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
f0  �a  �
�   $ ��  ��0  ��	�1  2�  �
�    I�  ��  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��1  ( 1  �1  =    ޴  �1  	�  .�  	�  /�  	�  0�  	�  2�  	w�  8f  	�  9-  	�  :�  	�_  ;�   	��  >�  	�  J�  	"�  R  	t�  S�   	�w  T�   	؜  Y�   	q�  [�  	Ƚ  ^  	�  _�   	�y  `�   	b�  c�   	+�  f�  	��  i�  	֘ l�   	�J  x�   	��  y�   	ks  �   	�  ��   	J�  ��   	�i  ��   	��  ��  	��  ��  	��  ��  	<� ��  	��  ��  	��  ��  	5�  ��  	<m  ��   	 K  ��   	�R  ��   	op  ��   	�m  ��   	D  ��   	X�  ��   	If  ��   	� ��   	��  ��  	�U  ��  	`  ��  	J�  ��  	��  ��  	� �G  �0  /4  =    	�  �4  �  K4  =    	� �;4  �  g4  =   	 	,�  �W4  	R�  �4  �  �  �4  =    	�u  ��4  	��  ��1  	�e  ��   �   �4  =   � 	(�  ��4  	�  ��   ��  G   �v  �    n�  �    4�  �    *b �    ��  �  �  ;5  ! 	R 05  �  R5  ! 	� G5  
K   $7  z  � �     & / 8 	; 
D M V _ h q z � q o z � � � � � � _ � o x �  � !�	 "  #1
 $� %< &( 'l
 (: )�	 *� +�
 ,� -V
 .# /� 0V 1� 2� 3� 4� 5a
 6� 7�
 8� 9� :D ;� <� =6 >f ?� @* Aa B C� D 
K   r�9  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	 V�   	�  �   	q  �9  �   	��  ��   	�\  ��  	�  ��9  �  	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  ��  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   C	�:  x E�   y F�   �{ H�:  (T	�:  `e V	   x W�  y X�  z Y�    	�  [�:  �a	�;  = c�   F�  d�  �~ eI  h�  fI  
t�  gI  �k hI  tag iI  �N  l
�   ��  o@0  ��  r
f0   iK  u�:  0��  x
�   XS�  {@0  `��  ~R   h��  ��   pu| ��<  x �}  X��<  v1 �R=   v2 �R=  dx ��  dy ��  �  �I  �k �I  tag �I  �W  �q  �o �X=  $��  �F=  4SX  �=  8d�  �=  @��  �
�   H��  �R   P �<  �;  �z �;  �	=  2�  ��   ]  ��  �h  �I  �N  �I  
�K  �I  >} �=   �<  �}  ��<  
K   �F=  ��   �  o�  ��   ��  �=  �:  �  h=  =    �u  ��;  �z ��-  8�	�=  v1 �R=   v2 �R=  82  ��  Mp �/  [�  ��=   �  ��=   SX  �=  (d�  �=  0 =  h=  A{ ��=  4	a>  %x �   %y 	�  %dx 
�  %dy �  �o a>  )�  �  0 �  w>  =   =    (} >  �  *�  &v  @2F?  @�  4F?   %x1 5�   %x2 6�   .]  8�  5]  9�  �� :�  ��  =�   �  @�   ��  C�  $�n  GL?  (9x  HL?  0�^  IL?  8 �=  I  >�  K�>  &�h  PR;@  s�  U;@   �H  V;@  %x1 X�   %x2 Y�   %gx \�  %gy ]�  %gz `�   %gzt a�  $�x  d�  (� f�  ,~�  i�  0t  k�  4.� l�   8�  pA@  @	�  r�   H _?  �>  �h  t_?  �	�@  �c  ��   �O  ��@  �x  �
�@   I  �@  =    �  �@  =    I�  �T@  �	�@  �  ��    �  ��@   �@  �  ��@  '��	�A    ��   �  �	�   t�  �	�   ��  �	�   /�  �	�   �  �	�  %top �	�A  (��  �	�  U(��  �	�  V(� �	�A  W(�  �	�  � �  �A  =   ? ��  ��@  	.L  &�A  �  	׮  )�A  	�  +�A  	�  ,�A  	�Q  .A@  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  76B  �   	��  86B  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�B  �@  	��  H�   	��  IR=  	��  K�   	a� LF?  	w�  N�   	P{ O=  	��  Q�   	��  R�B  t=  	��  T�   	�� UC  w>  	�}  W�   	u| X�=  	M�  Z�   	P�  [�=  	��  a�  	��  b�  	�  c�  	�p  e/  	�T  fzC  �0  	�a  j/  �   �C  =   � 	ը  l�C  /  �C  =   @ 	�p  m�C  	 �  p�  	p|  q/  	$Y  v�   	�K  y�   	g  {D  �A  	d�  |D  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   A@  �D  =   =   / 	��  E�D  A@  �D  =   / 	Ԁ  F�D  A@  �D  =   =    	7� G�D  	�R  I�   	��  JA@  	��  U�   	P�  \�  	��  ]�  	L�  ^�  	ߵ  _�  	�  a�  	@�  F?  	[�  �=  	 �  �=  	SX  =  	d�  =  	��  �   	_�   �   	��  "�  	��  %�  	'�  &�  	�]  (�  R?  �E  =   � 	�P  *�E  	ӯ  +F  R?  	|  -"F  A@  	��  ."F  	��  /"F  FF  VF  �   �    	��  L?  �   @F  	qY  "bF  	�  #bF  I  �F  =   ? 	��  %�F  	��  &�F  �  �F  =   � 	@Y  (�F  �  �F  =   ? 	V�  )�F  G@  �F  =    	�h  �F  	�  G  G@  	�  G@  	�f  !�F  	r�  "�F  	��  %L?  	��  &L?  	׆  '�  	��  (�  	�  *�  	��  +�  	�   A@  	��   �   	�_   �   	�_   �   	b   �  	t   �  	j�   "�  	�   :�   	��   ;�   	��   <�   	�W   >A@  	hn   @�  	U~   A�  	�   B�  	 �   C�  	%�   F�  	�u   H�  	z   I�  	ʓ  !C	  �  vH  =    	��  !bfH  �   �H  =    	��  !c�H  	0K  !d�   	?�  !e�   !�	�H  x !��   y !��  dx !��  dy !��   ��  !��H  !�I  �p !�
@0  ��  !�
�=   !�	KI  {q !��   ��  !��  d !�	�H   t�  !�I  KI  gI  =   � 	r !�WI  	�T  !�I  KI  	l�  !��  	�  !��  	?k  !��  	�d  !��  	2~ !��H  	��  !��  	��  !��  	k�  !��  	Z�  !��=  �=  J  =    	�v  !��I  	�v  !��   	"�  !�@0   �  !�   �U  !L?   ��  !L?   t�  !�    �  !	�    .Y  !
�   7Y  !�   �h  !�J  @0   *� !f0   <i  !f0  	G  "�  	��  "�   
K   "��J  )top  �G  �  �]  "��J   "�	=K  ��  "��=   ��  "��J  O{  "�
�   ��  "�
�   iK  "�=K   �:  ��  "��J  CK  _K  =    	��  "�OK  "K   "�K  )up  �  �F  �S   FT  "
kK  "K   "�K  ��   �x  H�  ��  �H   ��  "�K  H"	�L  `e "	   >} "=  L� "�   %low "�  $+� " �  (�Z "!
�   ,r� ""
�   0�f  "#�K  4�f  "$�K  8��  "%�  <%tag "&
�   @*� "'�K  D �w ")�K  �L  �L  =    �L   �  "2�L  "K   "��L  ��   �s  z�  ��  �T  ܭ   gY  "��L  H"�	�M  `e "�	   *� "��L  >} "�=   �W  "��  (�}  "��  ,L� "��  0��  "��  4��  "�
�   8%tag "�
�   <��  "�
�   @  w "��L  �M  �M  =    �M   j�  "�M  =� #�M  ��  #.N  ^�  #2�N   }�  #7�  �� #;K    #	7N  r� # LN   .� #$]N  O� #)�N   *FN  FN  �    �M  7N  ]N  FN   RN  *1   �N  FN  K   R   1    cN  ��  #,N  �N  oS  $'�N  dS  ($)O  � $+
a   � $,FN  @�  $-
�   >z $.
�   �  $/R   �H  $3O    �N  	�� $7O  	�� $8K   
K   %"dO  ��  WH  �~  �O  �m  ��   �  ��  ��  	 B	�O  �@ EI   �� H@0  t K	�    ]� MdO  + Q�O  	x%f     �O  ,�2  V	t�e     ,�2  Z	p�e     +@� ^�   	t%f     +8� b�  	p%f     +ƞ f#P  	h%f     �  ,�9  j	l�e     -מ �$�A     Z       ��P  .=�A     �Y  .B�A     �Y  .R�A     �Y  .a�A     �Y   /�� �	�  �A            ��P  0$�A     
Z   -L Y~�A     �       ��Q  1C� Y�   �I �I 1? Y&�   (J J 2� [#P  �J �J 3��  \
9  �W2t ]R   �J �J 4��A     Z  bQ  5U	�B      .��A     ;P  4��A     "Z  �Q  5U�W5T95Q	'�B      4��A     .Z  �Q  5U�W 4�A     :Z  �Q  5T1 .�A     FZ  .%�A     RZ  63�A     ^Z  5Tv   -n T��A            �FR  1Ҟ T�   �J �J 7��A     �P  5U�U5T0  -E\ Fh�A            ��R  1Ml  F�   =K 7K 6~�A     Z  5U	��B     5Ts   -�X ;J�A            �S  1Ml  ;�   �K �K 4`�A     Z  �R  5U	��B     5Ts  7h�A     jZ  5U�U  -� ���A     �       �
T  1b� �@0  �K �K 2� ��   IL GL 2�k ��   vL lL 3Ml  ��   �H8sep ��   �L9sfx �I  �L �L 9c ��O  M M .��A     vZ  .��A     �Z  4�A     %V  �S  5U| 5Q�H5R�L .,�A     �Z  .5�A     SX   -& �[�A     &       �7T  .t�A     �Y   -$" �5�A     &       �dT  .N�A     �Z   -� �i�A     �      �%V  1g� �R   9M 3M 1k� �'�   �M �M :sfx �I  2�� �@0  �M �M 9rc �	�   +N )N 8sep �	�   �H2�k �	�   PN NN 3Ml  �	�   �L;W  D�A     �  ��U  <2W  =%W  uN sN >�  ??W  �N �N ?LW  )O 'O 4o�A     SX  {U  5U}  6��A     SX  5U}    4��A     Z  �U  5U	��B     5Ts  4 �A     %V  �U  5T| 5Q�L5R�H 4D�A     XW  �U  5U|  4
�A     �Z  
V  5Us  6'�A     �Z  5Us 5T}   @N� C�   &�A           �W  1b� C(@0  RO LO 1m�  C:@0  �O �O Avol D%6B  �O �O Asep D/6B  3P -P 2L� F�  �P P 9adx G�  �P �P 9ady H�  4Q 2Q 2Mp I/  [Q WQ .��A     �Z  6��A     �Z  5UHB$  B� �   XW  C�� !@0  C�@ 4I  D�k 	�   :c �O   E(t �:�A     /       ��W  F�� �@0  �Q �Q G�k �	�   �Q �Q 0`�A     SX   E�| �A�A     �       �CX  G�k �	�   ?R 7R GX� �	�   �R �R H��A     -       X  +� �CX  �L 4h�A     SX  /X  5Us  7��A     �P  5T1  �   SX  =    I|� ���A     8       ��X  F�k ��   �R �R Ji �	�   S S Jc ��O  =S ;S .�A     �Z  .�A     �Z   E�� ���A            ��X  .��A     �Z  0��A     �Z   E�
 r��A     �       ��Y  F�J  r�   fS `S F��  r �   �S �S Ji t	�   
T T 4��A     �Z  mY  5Tm 4��A     FR  �Y  5Uv  4��A     �R  �Y  5Us  4��A     [  �Y  5T15Q0 7�A     [  5U	��A     5T1  K�? �? �K�> �> �K.? .? �K} } $I	K�> �> �	K��  ��  &7KG�  G�  '/K�{ �{ $=K� � $BK�} �} $?K�? �? �K#? #? �Kb> b> �K?? ?? �K
? 
? �	K�@ �@ �KM? M? �K�@ �@ �K�? �? �KEf Ef xKd  d  "	K7> 7> �K@ @ �KY? Y? �K�= �= �K� � %6K  &A 	   ��  S#  � �*  ��A     )       5� �  ,	  0t  D   e2    �  �0  }  int ^&  ��  8   ڵ  Ru   �   t�   g   �   �   �   1   �' �   ��  1�   ]  4�   	�   �   �   1   � �   Zy  8�   �     
1   
1   � �   ��  ;  Ʃ  QR      ,  B  1     1  �  WB  �   @	��C     �   E	��B     �   I	x�e     G  K	��B       Q	��B     �� )g   ��A     )       �num )R   XT TT den )-R   �T �T ans +R   �T �T   �   t�  S#  �� �*  ��A     s      2� ��  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  �� �  0t  ;  e2    �0  }  ��  /  
K   J�  D   �C  
D  ���� �C  Nc  ڵ  RW  �  	��  ��   	�\  ��  	�  �(  	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  ��  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   (	�  ��  P      P  Vd  !P  �  "P  �� #�   �   �  =    � %Y  (	�  � *�   �� +�   � ,�  G /�  �     =    	N�  	%�  	��  	'�  P� 	,0  6  �  O  O  �   �    �  =� 
a  ��  
.�  ^�  
2#   }�  
7�  �� 
;K    
	�  r� 
 �   .� 
$�  O� 
)   �  �  �    U  �  �  �   �  1     �  K   R   1    �  ��  
,�    oS  '5  dS  ()�  � +
�   � ,�  @�  -
�   >z .
�   �  /R   �H  3�    �   �  =    )  	�� 7�  	�� 8K   
K   "  ��  WH  �~  �O  �m  ��   �  ��  ��  	   3	�%f     {� 6�  	�%f     �� :�  	�%f       <	�i     � @$  	�%f     �n	c  � p�    �  q�   � r�   �� s�   F� uB  >� vB  f� wB  ,� xB  
-� zB  ܠ {B  @� }c  $� �   @g� ��   A� �B  B"� �B  Dt� �s  F"8 �;  � ;  s  =   / �   �  =   9 a� �j  �	 N��A     �      �f	  L� N�   �T �T 1� P�   �� Q	�   vU rU :� Q�   �U �U red Q�   V �U ǡ Q$�   gV aV �� Q+�   �V �V ͡ Q2�   /W )W 2� R	�   zW xW 8� R�   �W �W C� S	�   �W �W �� T	�   X X ԡ U	�   /X +X ��A     ?  �  UwTwQw ��A     ?     UUTUQU ��A     ?  "  U�T0Q0  B     ?  C  U0T0Q0  B     ?  f  U�T�Q0 2 B     ?  �  U�T�Q� � B     �  �  U�T?Qq Rr Xx  � B     e  �  U�T?QxR9X  � B     �  	  U�TCQq Rr  B     �  3	  U�TCQq   4B     �  !YB     o  U�T@Qq Rr   3 6�A     v       ��
  %� �   kX eX i 	�   �X �X "Ġ 
�
  �P#ext �   
x�C     �[�A     K  
  Uw T@Qv Rs X	x�C      c�A     W  #
  Uw  z�A     c  B
  U	|�C      ��A     o  f
  U	�RB     T8 $��A     �
  Uw Q
@R�  �   �
  =    � �)�A           ��  ��  ��   �X �X "8 �)�  RY DY ��  ��   
Z Z   �"�   \Z VZ @� ��  �Z �Z i �
�   W[ I[ �� �
�   �[ �[ pcx ��  %\ \ ��  ��  �\ n\ c�A     {  �  U~ 1$#�T1Q0  �A     �  �  Uv Ts  %6�A     �   �  &� e�A            �w� ^�A            �  '�< ^�  U &4 U�A            �y� M��A            �e  (raw M�  �] �]  �� @��A     :       �o  (x @�   �] �] (y @�   ^ ^ (w @"�   W^ Q^ (h @)�   �^ �^ )c @0�   X��A     �    Uz Ty Qq Rx  ��A     �  *  Uz Ty { "1 ��A     o  N  Uz Ty Qq  !��A     o  Uz �Q"1Ty   �� 2��A     ,       ��  (x 2�   �^ �^ (y 2 �   _ _ )h 2'�   Q)c 2.�   Rbuf 4�  __ W_ y1 5	�   �_ �_  W  � %t�A     %       ��  )x %�   U(y %!�   ` ` )w %(�   Q)c %/�   Rbuf '�  U` M` x1 (	�   �` �`  ̠ :�A     :       �@  (x �   a a (y !�   Ta Pa )w (�   Q)h /�   R)c 6�   Xbuf �  �a �a K� �  �a �a x1 	�   Pb Jb y1 �   �b �b  & ���A     �       �   (x ��   �b �b (y ��   0c (c ��  �$�   �c �c   �/�   �c �c (src �=�  #d d `5 ��  �d d ��A     c  �  U	h�C      $�A       U~ T�TQv R}   �� ���A            �`  $��A     o  U	a�C     T1  �� �}�A            ��  $��A     o  U	Y�C     T1  � ���A     �       ��  (x ��   �d �d (y �%�   Ue Oe .� �1O  �e �e r� �	�   �e �e col ��   cf [f � ��  �f �f � ��  �f �f `5 ��  tg lg m�  ��  �g �g �� ��  ih ]h M9 ��  i �h w �	�   ti ri $��A     c  U	A�C       �  �� z��A     �       ��  (x z�   �i �i (y z"�   j  j .� z/O  Xj Rj r� |	�   �j �j col |�   �j �j � }�  2k 0k � ~�  _k Uk `5 ~�  �k �k m�  ~�  4l ,l w 	�   �l �l $��A     c  U	,�C       � I��A     �       ��  (x I�   �l �l (y I �   m m .� I-O  |m rm r� K	�   �m �m col K�   n n � L�  in en � M�  �n �n `5 M�  �n �n m�  M�  Mo Go w N	�   �o �o *7�A     Uv T| Qs   k� �A     �       ��  (x �   �o �o (y �   Ap ;p .� ,O  �p �p r� 	�   �p �p col �   q q � �  mq kq � �  �q �q `5 �  r r m�  �  or gr w 	�   �r �r $a�A     c  U	�C       � �A            �k  (x �   �r �r (y #�   5s 1s .� /O  rs ns !�A     �  U�UT�TQ�Q  + �"�A     �       ��  ,x ��   �s �s ,y �$�   t �s -.� �0O  nt dt .r� �	�   �t �t /col �	�   Nu Hu .� ��  �u �u .� ��  �u �u .`5 ��  7v /v .m�  ��  �v �v /w �	�   +w )w 0W�A     k  Uv T| Qs  ��A     c  �  U	�C      $��A       U|   +y�  � �A           ��  ,x ��   Tw Nw ,y ��   �w �w -.� �)O  x x .r� �	�   �x �x /col �	�   �x �x .� ��  ?y =y .� ��  jy by .`5 ��  �y �y .m�  ��  Yz Qz /w �	�   �z �z 0^�A     �  Uv T| Qs  ��A     c  �  U	��C     T| Qs  $��A       U|   +�� ��A            �  1ڈ �.$  U +1� U@�A     �       �  -�� U�   �z �z -¡ U�   I{ C{ -m�  U+�  �{ �{ -��  V�   �{ �{ -  V �   '| #| -/� W�   c| ]| 15� W �   � /src Y�  �| �| .`5 Z�  } } ��A     c  �  U	��C      $��A       U Ts Q| R}   2��  EY  3x E�   3y E�   4��  E#�   4  E.�    5  ��A     K       �?  6,  C} ;} 66  �} �} 6@  &~ ~ 6L  �~ �~ 7  @  6L  �~ �~ 6@  B > 86  6,  � { $�A     �    U	�i     Ts Qv  !?�A     �  U	�i     T	�U�Q"1Q	�T�R"1   9T� T� i9G�  G�  /9$�  $�   	9��  ��  79��  ��  C9� � 69�. �. 	9� � 7	9�L �L ) 1n   ��  S#  A� �*  hB     �      j� ��  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  
K   "f  ��  WH  �~  �O  �m  ��   �  ��  ��  	 0t  r  e2    �0  }  ��  f  
K   J�  D   �C  
D  ���� �C  N�  ڵ  R�  �  	"|  *�  	��  +�  	I�  ,�  	�a  -�  	 	�  ��  	"�   E�  	#�  e% 	$�  u  	%
�  �8 	&
�  ��  	)
�  /b  	-
�  ��  	.	�   a  	2
�  �T  	3
�   Mx 	4  
K   
!�  �p   �  ��  S�  ��   �F  
'�  
*	'  *� 
,�   "G  
C	�   (G  
C�   �]  
C�   :G  
C�    �U  
D�  
K   
K�  � � ^�  �� e  2 8� ��  �  _�  �   �  
K   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  
K   /  ��   [r  �4 #�  �   �X  5�  
K   :~  7g   G�  Dg  Qg  ^g  %�  h  �l  �E  ��  	��  
��  ��  ��   ;�  K  
�   P�  =_  ��   R�  N�  ��  ��   �p  W�  =� �  ��  .
  ^�  2�   }�  7�  �� ;K    	;  r�  P   .� $a  O� )�   J  J  �    �  ;  a  J   V  1   �  J  K   R   1    g  ��  ,
  �  �  oS  '�  dS  ()  � +
   � ,J  @�  -
�   >z .
�   �  /R   �H  3    �     =    �  	�� 7  	�� 8K   
K   3`  ��   ({  ��  ğ   F]  89  
K   Y�  ��   �c  |  ��  l  ��  �   
K   k�  _   �m  ��  }  �  �f  TO  #�  �  oT  	B�  
 {�  {�  
K   �5  &�   �  º  GY  �f  ��   v�  �  
K   �z  GQ   ϼ  �  �_  X  &�  �b   	� M�   	5 N�   t�   �   �  �  �  =   �' �  	��  1�  	]  4�  �  �  �  =   � �  	Zy  8�  �    =   =   � �  	��  ;  Ʃ  QK      ,  B  =     1  	�  WB  �p  #_  e  l   S�  $x  ~  �  R    T}  %�  �  �  R   R    '	�  acv )S  ��  *l  ��  +�   �y -�  �Y  6�  ��  :&	  s�  <&	   �H  =&	  xz  >�   �  x @�  �  H	  =    y  X	  =    
�	�	  x ��   y ��  Mp ��  *� ��  ޽  ��   ~x �X	  
K   �  @�   9�  �E  C�  �p  0�  ��  �r  zr  �U  	�U  
�O  	�   �  ��  ��  A�  �  /�  8�  1�  ��  �U  �  �  �  �  ;�  I�  �  	i  ��  7�   i�  !�s  "$�  #��  $��  %��  &ٗ  'v�  (a�  )+�  *Rr  +Ϝ  ,p�  -Զ  .�p  /�b  0ҟ  1��  2�  3�U  4A  5�  6�  7#�  8�  9��  :��  ;�  <
�  =Tc  >�  ?��  @��  A�j  B�]  C�  D��  E�  F��  GK�  H��  I.�  JL�  K0x  L x  M��  N�  O��  P�T  Q��  R��  SA�  T�  U��  V��  W�F  X=o  Y�E  Z��  [	�  \{s  ](^  ^�  _�P  `R�  a[�  b��  c��  dI�  ed�  f�P  g�P  h�P  i�P  j��  k�]  lS�  m�]  n�]  o��  pQ  q�]  r��  s��  t��  u��  vm�  w�]  x8  yJ�  zA�  {��  |z�  }�  ~د  �  ��  ��  ���  ��  ��  ��  ��Y  ��  � �  ��X  � �  ��	  
K   ��&  �Q   
�  �e  R�  ��  ��  ��  �  �  �  	�X  
8�  h�  ��  *�  ��  ��  ��  	Q  V\  ��  ��  ��  ��  ��  ��  ��  ��  ś  ͛  �g  �g  4i   Tw  !|  "�  #��  $��  %��  &��  '��  (��  )��  *��  +H  ,�G  -{�  .�  /��  0��  1%�  2��  3&�  4/�  58�  6c�  7q�  8�J  9z  :�K  ;�d  <�d  =�d  >�P  ?��  @�P  A��  BX  C�J  D��  E.�  F��  G��  H�  I�R  J�H  K�X  L�J  M�J  N^`  Om`  P  Q��  Rd�  S&d  T-d  U4d  V;d  W!�  X-�  Yc�  Z�o  [�o  \��  ]wl  ^��  _��  `L�  aU�  bad  ckd  dud  e�y  f�y  gQ�  h[�  ie�  j]  k_�  l8�  m�  n�  o�  p��  q_  rܸ  s��  t��  ut�  v�  w��  x��  y��  z��  {<�  |F�  }P�  ~��  ��  ���  ��d  �ݶ  ��  �ڬ  ��  ��  ��  ���  ��  �
�  ��  �,�  �u  ��h  ��h  ���  ��  ��  ��  ���  ���  ���  ���  ���  �Y  �Y  �k�  �A�  �Wf  �cf  �of  �{f  ��f  ��f  �f�  ��m  ��m  � n  �n  �n  �'n  �4n  �An  �Nn  ���  ��  ��{  ��{  ��{  ��{  ��{  ��{  ��{  � |  �k�  �w�  ���  ���  ��  �D�  �P�  �\�  �|a  �s�  �)�  �6�  �C�  �ӿ  �P�  ��  �k�  ���  ���  ��  �(�  �6�  �D�  �(i  ���  �&a  �2a  ���  �>a  ���  ���  �Qa  ���  ��  ��  ���  �w�  ���  ���  ���  �  �Ύ  �ڎ  �&U  �3U  �@U  �MU  �ZU  �gU  �tU  ��U  ��U  �P�  �^�  �l�  �z�  ���  �'�  ��  ���  ���  ��~  ��~  ��~  ��~  ��~  �׈  ��~  �7�  �D�  �Q�  ��  �*�   6�  B�  �^  X�  d�  p�  |�  �  Z�  	y�  
��  ��  ��  8b  ��  G  ų  ѳ  ݳ  �  I|  @G  d|  ĵ  l  l  �  $l  ,l  4l  <l  X�   Tl  !��  "��  #��  $��  %��  &��  '��  (��  )�  *�  +)�  ,2�  -;�  .D�  /M�  0V�  1_�  2h�  3q�  4z�  5��  6��  7�  8=�  9�  :!�  ;*�  <��  =�  >i�  ?X�  @��  A�  Bя  Cݏ  D�  E��  F�  G�  H�  I%�  J1�  K��  L��  M��  Nz}  O��  P�}  Q�}  R�e  S�e  Tɇ  Uև  V�F  WSx  X'�  YM�  Z3�  [?�  \b  ]T�  ^v�  _��  `��  a��  b��  c��  dy  ey  f�_  g�_  h�r  i��  j	�  kG�  lS�  m.G  n_�  ok�  pw�  q=|  rVG  s��  tj�  uw�  v+  wR�  x^�  yj�  zv�  {��  |��  }��  ~��  ��  ��  �=f  ��h  �=~  �I~  ���  ���  �~~  ���  �A�  �M�  �?�  ��  ���  �
�  ��  �&�  �4�  �B�  �P�  �^�  ���  �y�  �[�  �g�  �s�  ��  ���  ���  ���  ���  ���  ���  ���  ���  �^�  �}b  ���  �
�  ��  �"�  �.�  �:�  �q�  ���  ���  ���  ���  �Ԗ  ��  ��M  ��M  �N  �?�  �N  �-N  �;N  �L  ���  �q�  �}�  ���  ���  ���  ���  ���  ���  �zS  ��S  ��S  ���  ��i  �0m  ��`  ��`  ��`  ��`  �˞  �؞  ��  ��  ���  ���  ���  ��  ���  �
�  ��  �&�  �4�  ��h  �{w  �K  �K  ���  �r�  �9K  �EK  �QK  �]K  �Fo  �Ro  �^o  �u�  ��  �d{  �p{  �|{  ��{  ��{  ��{  ���  �ǥ  �ե  ��  ��  ���  �J  �^�  �߄  ��  ���  ���  �s�  ���  �M�  �Y�  �e�   �  q�  }�  ��  ��  ��  ��  S�  rj  	`�  
j�  ��  ��  >�  nr  ��   �  ,�  8�  D�  P�  \�  h�  t�  ��  ��  ��  &e  S�  )�  5�  A�   /q  !M�  "Y�  #e�  $S  %S  &S  ',S  (:S  )HS  *VS  +͗  ,��  -�z  .�z  /�z  0�z  1�z  2�z  3{  4{  5R�  6^�  7j�  8��  9�  :H�  ;T�  <`�  =l�  >x�  ?��  @��  A�E  B�E  C�E  D�E  E�E  F�E  G	F  H�}  IԷ  J�  K��  LS�  Mf�  Nt�  Og�  P��  QT�  R)�  S6�  TC�  UP�  VIN  WVN  X�a  Y�e  Zv�  [��  \�  ]+�  ^7�  _��  `K�  aW�  bc�  cN�  d[�  eh�  f��  g�Q  h�Q  ikg  j�  kK�  lCu  mOu  n[u  ogu  pfj  qsu  ru  s�u  t�u  u��  v��  wnG  xm�  y�x  z��  {��  |��  }��  ~�  �  ��  �)�  �5�  ���  �ʊ  �׊  �P  �P  �P  ��d  ���  �l  �k]  ��  �3�  �S�  �_�  �w�  ��  �q  �q  �!q  ���  �;q  �v�  �`q  ��  ���  �W�  ���  ��  ���  ���  �5�  ���  ��  �k�  ��  �(�  �5�  �B�  �O�  �\�  �H�  �U�  �b�  �o�  �|�  ���  �jQ  ��  ��  �'�  �4�  �A�  �N�  �[�  �h�  �u�  �mw  �Y�  ���  ���  ���  ���  ���  ���  ���  ���  ��w  ���  ��}  �:�  �=P  �IP  �UP  �aP  �mP  �yP  ���  ���  ���  � �  ��  ��  �d�  ���  �]m  �im  �um  ���  ��m  ��m  ��m  ��m  �*�  �6�  �B�  �N�  �Z�  �f�  �s�  ���  ��  ��  ��  �(�  �4�  ���  �Π  ���  ���  �nq  �{q  ��q  ��q  ��q  ���  ���  ���  ���  ���  ��  ���  ���  ���  ���  ���   ȕ  ԕ  ��  �  ��  Eb  Rb  �  wQ  	��  
�P  D�  ��  ��  ��  da  �R  bG  ]�  f�  o�  �  ��  �  ��  ��  ��  ��  ǀ  3�  ��  �   �  !zT  "!H  #�T  $(K  %��  &��  '�  (OY  )WY  *_Y  +�r  ,t�  -|�  .��  /lb  0��  1��  2fr  3��  4Ĩ  5B�  6�t  7�t  8��  9��  :��  ;��  <Jr  =4�  >ܣ  ?��  @1�  A[O  B��  C�N  DI�  E��  FI�  G�T  H�  I��  J�o  K�o  L�o  M�o  N�o  O��  P`�  Qh�  Rj�  S��  T��  U�G  VZ�  W�G  X��  Y$�  Z,�  [4�  \|�  ]�J  ^�  _�  `�~  a#�  b+�  cmH  d%Q  e!h  f�  g��  h��  i�  j��  k4�  l>t  m��  n�w  oB�  pj�  q��  r͖  s��  tC�  u��  v�y  w�  xN`  yD�  zT�  {�U  |*�  }d  ~R�  {�  ��o  ��  ���  �V  �m}  ��X  ��X  ��X  ��  �{Y  ��  ��]  ���  �҅  ���  �^�  �Ĝ  ��j  �۾  ��|  ��X  ���  ���  ���  ��  ���  ���  � �  ���  ���  �f�  �s�  ���  �3�  ���  ��  ��  �9�  ��  ���  ��  �	O  ���  �>�  �'�  ���  ��N  ��N  ��N  ���  �s�  ���  ���  ���  ��y  �z�  ��G  ���  �+�  �Jd  �ҽ  ���  ���  ��r  ��  ��  ���  ���  ���  ���  �ߤ  � ��  u  (x		'   �u z�    � {	�    s |	�    � ~�   N�  �&   ��  �	�    ��  �	�     J]  ��&  	'  ''  =   � !�^  �'  �   ?'  " !�  �4'  #K   ��*  q�   �R  �z  ��  Bd  g�  LG  g�  p�  ��  	*�  
�z  =�  �Q  jv  �a  V�  Z�  3�  ��  ��  ��  �f  ��  ��  ��  �t  ��  i�  �s  �r  X�  ��   o�  !�  "�q  #gh  $��  %�l  &��  ',�  (��  )��  *�  +�  ,&�  -/�  .8�  /A�  0J�  1�\  2�\  3�\  4�j  5�f  6�j  7]a  8�f  9Ja  :�j  ;�f  <k  =l�  >��  ?!k  @+k  A5k  B�l  C�l  D<h  E�l  F�l  G�l  H��  Im  Jm  Km  L�z  M'�  N&m  O�n  P��  Q�n  R�n  S o  T
o  Uo  V�  W)o  X3o  Yep  Z�s  [}p  \�p  ]��  ^��  _�p  `��  a�s  b�p  c�q  dq�  e�q  fr  gr  hr  i"r  j,r  k6r  l@r  m�r  n�r  o{  ps  qs  r s  s*s  t4s  u>s  vHs  wEt  x��  yOt  zYt  {ct  |mt  }wt  ~  �t  ��t  ���  � v  �*v  �4v  �>v  �Hv  �Rv  �th  � o  L'  \	�+   �Y  	�     *O  	�    ��  	�    �  	�    b�  	�    ��  	�    �  	�    +�  	�    Zp  	�     o�   	�   $ m�  !	�   ( 4�  "	�   , �  #	�   0 �  $	�   4 ��  %	�   8 L� &	�   < ��  '	�   @   (	�   D ��  )	�   H \q *	�   L z�  +	�   P �  ,	�   T /�  -	�   X ʤ  /�*  �+  ,  =   � !��  1�+  �]  ���-  `e �,	   x ��  y ��  z ��   ��  ��-  (cN  ��-  0Mp �   8�u ��  <� ��   @�H  ��-  Hr�  ��-  P��  �-.  X��  ��  `m�  ��  d��  ��  h  ��  l3F  ��  p8F  ��  t=F  ��  x��  ��   |*� ��*  �y� �3.  �s ��   ��� �9.  ��  ��   ��  ��   �ʺ  ��   ��l  ��   �  �  �-  � ��  �   � ��  	�   � �R  0  � f�  �   � I}  �	  � ��  �-  � ,  Gx  �-.  >} ��3   �}  ��  �|  ��  
 �-  �+  	'  $d  HN0  mo P�2   ��  Q�9  cmd R�  �  W�  (_  Y�   #_  [�  $bob ]�  (�  a�   ,�[  b�   0sb  d�   4d]  g�9  8�W  h�9  P��  i�  h�� l�2  l�N  m�  |E�  p�  ��W  r�9  �~�  s�2  �*� t�2  ��� w�   ���  x�   �X�  |�   ��e  �   ���  ��   �g  ��   ��u  ��   �|G ��   �Q  ��   ��  ��   �o�  ��2  �%�R  ��    %��  ��   %�  ��   %h  ��9  %I�  ��  @ ?.  �z ,  	��  ��   	�\  ��  	�  �P0  �  	��  ��   	��  ��   	2�  ��  	��  ��   	Ɇ  ��  	��  ��   	��  ��   	�h  ��   	rK  ��   	l�  ��   	]�  ��   	��  ��   (	21  ��  �      �  Vd  !�  �  "�  �� #21   �   B1  =    � %�0  C	n1  x E�   y F�   �{ HN1  (T	�1  `e V,	   x W�  y X�  z Y�    	�  [z1  �a	�2  = c�   F�  d�  �~ e�  h�  f�  
t�  g�  �k h�  tag i�  �N  l
�   ��  o�2  ��  r
�2   iK  u�1  0��  x
�   XS�  {�2  `��  ~R   h��  ��   pu| �n3  x 0  �   �2  =    �}  X�n3  v1 �#4   v2 �#4  dx ��  dy ��  �  ��  �k ��  tag ��  �W  �8	  �o �)4  $��  �4  4SX  ��3  8d�  ��3  @��  �
�   H��  �R   P t3  �2  �z ��1  �	�3  2�  ��   ]  ��  �h  ��  �N  ��  
�K  ��  >} ��3   z3  �}  ��3  
K   �4  ��   �  o�  ��   ��  ��3  n1  �  94  =    �u  ��2  �z ��-  8�	�4  v1 �#4   v2 �#4  82  ��  Mp �   [�  ��4   �  ��4   SX  ��3  (d�  ��3  0 �3  94  A{ �Q4  4	25  &x �   &y 	�  &dx 
�  &dy �   �o 25   )�  H	  0 �  H5  =   =    (} �4  �  *�  'v  @26   @�  46   &x1 5�   &x2 6�    .]  8�   5]  9�   �� :�   ��  =�    �  @�    ��  C�  $ �n  G6  ( 9x  H6  0 �^  I6  8 �4  �  >�  Kb5  '�h  PR7   s�  U7    �H  V7  &x1 X�   &x2 Y�   &gx \�  &gy ]�  &gz `�   &gzt a�  $ �x  d�  ( � f�  , ~�  i�  0 t  k�  4 .� l�   8 �  p7  @ 	�  r�   H 06  U5  �h  t06  �	Z7   �c  ��    �O  �Z7   �x  �
j7   �  j7  =    �  z7  =    I�  �%7  �	�7   �  ��     �  ��7   z7  �  ��7  (��	k8     ��    �  �	�    t�  �	�    ��  �	�    /�  �	�    �  �	�  &top �	k8  )��  �	�  U)��  �	�  V)� �	k8  W)�  �	�  � �  |8  =   ? ��  ��7  	�8  ~�  5   �S  
�   ��   
�     !
�   �g  "
�   �^  #
�    ��  %�8  �8  �8  =    	S�  '�8  
K   7*9  {�   U�  ~�   >	f9  �� @9.   s A
�   sx B�  sy C�   Nz E*9  
K   1�9  ��   ��  ��   �y  9r9  �   �9  =    �  �9  =    �  �9  =    f9  �9  =    hy �?.  (�	O:  in ��   d  �
�   �x  �
�   D  �
�   5O  �
�   �� �
�2  �a  �
�   $ ��  ��9  ��	�:  2�  �
�    I�  ��  r�  �
�   �H  �
�   *F  �
�   ��  �
�   	�  �
�   ѵ  �
�   ��  �
�    F� �
�   $�  ��:  ( O:  ;  =    ޴  �[:  	.L  &;  �  	׮  );  	�  +;  	�  ,;  	�Q  .7  	��  0�   	��  1�   	(_  2�   	դ  4�   	�j  7�;  �   	��  8�;  	@�  <�   	�O  =�   	(g  >�   	�^  E�   	�u F�;  �7  	��  H�   	��  I#4  	��  K�   	a� L6  	w�  N�   	P{ O�3  	��  Q�   	��  RB<  E4  	��  T�   	�� U`<  H5  	�}  W�   	u| X�4  	M�  Z�   	P�  [�4  	��  a�  	��  b�  	�  c�  	�p  e   	�T  f�<  �9  	�a  j   �   �<  =   � 	ը  l�<     =  =   @ 	�p  m=  	 �  p�  	p|  q   	$Y  v�   	�K  y�   	g  {Z=  |8  	d�  |Z=  	��   �  		�  !�  	�3 #�   	_  $�   	-�  (�   	�f  )�   	�G  +�  	`�  ,�  	A�  -�  	��  /�   	��  1�   	P�  2�   7  >  =   =   / 	��  E�=  7  .>  =   / 	Ԁ  F>  7  P>  =   =    	7� G:>  	�R  I�   	��  J7  	��  U�   	P�  \�  	��  ]�  	L�  ^�  	ߵ  _�  	�  a�  	@�  6  	[�  �4  	 �  �4  	SX  �3  	d�  �3  	��  �   	_�   �   	��  "�  	��  %�  	'�  &�  	�]  (�  #6  P?  =   � 	�P  *@?  	ӯ  +h?  #6  	|  -z?  7  	��  .z?  	��  /z?  �?  �?  �   �    	��  6  �   �?  	qY  "�?  	�  #�?  �  �?  =   ? 	��  %�?  	��  &�?  �  @  =   � 	@Y  (@  �  4@  =   ? 	V�  )#@  7  P@  =    	�h   @@  	�   h@  7  	�   7  	�f   !�?  	r�   "�?  	��   %6  	��   &6  	׆   '�  	��   (�  	�   *�  	��   +�  	�  !7  	��  !�   	�_  !�   	�_  !�   	b  !�  	t  !�  	j�  !"�  	�  !:�   	��  !;�   	��  !<�   	�W  !>7  	hn  !@�  	U~  !A�  	�  !B�  	 �  !C�  	%�  !F�  	�u  !H�  	z  !I�  ) "�A  J @"NB  � ""�    � "'
NB  �� "*	�   
 "-^B  �9 "0	�    Ml  "3	�   $	
 "8	�   (C� ";	�   ,� "?	�   0� "BR   8 �   ^B  =    �A   "H	�B  � "K�    C� "N	�   "8 "QR   t "TR    . "VdB  	: "��   	3 "��   	� "��   	� "��   	O "��   	�
 "��   �A  C  " 	R #�B  �B  C  " 	� #C  
K   #$�D  z  � �     & / 8 	; 
D M V _ h q z � q o z � � � � � � _ � o x �  � !�	 "  #1
 $� %< &( 'l
 (: )�	 *� +�
 ,� -V
 .# /� 0V 1� 2� 3� 4� 5a
 6� 7�
 8� 9� :D ;� <� =6 >f ?� @* Aa B C� D 
K   #rtG  �  6  -   A D � � 	2 
� � � q � � � _ $ �  + � � v � � � x � ` �  Z !� "� #� $� %� &� '� (� ) *� +� ,� -x .� /� 0P 1� 2� 3  4� 5
 6� 7| 86 9� :� ;� <� =[ >j ?' @� A BO C� D� E" F� Gc H` I� JF K L� MA N< O� Pn Qt R� SL T� U� V� WU X0 Y� Z [� \� ]{ ^ _� ` a. bJ ci d e: f  g� hf i� j� k lK m 	 $V�   �  	��  %M�  	(h  %N�   	l�  %N�   	�  &.�  	�  &/�  	�  &0�  	�  &2�  	w�  &8  	�  &9�  	�  &:~  	�_  &;�   	��  &>�  	�  &J�  	"�  &R�  	t�  &S�   	�w  &T�   	؜  &Y�   	q�  &[�  	Ƚ  &^�  	�  &_�   	�y  &`�   	b�  &c�   	+�  &f�  	��  &i�  	֘ &l�   	�J  &x�   	��  &y�   	ks  &�   	�  &��   	J�  &��   	�i  &��   	��  &��  	��  &��  	��  &��  	<� &��  	��  &��  	��  &��  	5�  &��  	<m  &��   	 K  &��   	�R  &��   	op  &��   	�m  &��   	D  &��   	X�  &��   	If  &��   	� &��   	��  &��  	�U  &��  	`  &��  	J�  &��  	��  &��  	� &�`  �9  J  =    	�  &�J  �  .J  =    	� &�J  �	  JJ  =   	 	,�  &�:J  	R�  &�bJ  �	  �	  xJ  =    	�u  &�hJ  	��  &�;  	�e  &��   �   �J  =   � 	(�  &��J  	�  &��  !��  &`  !�v  &�   !n�  &�   !4�  &�   !*b &�   !��  &�G  	N�  '%�2  	��  ''�  B1  
�   (RK  6� B�  ٦  � (!1K  
K   nK  ��  �� �  ޣ s^K  u	�K  x w
�    y x
�    "�  z�K  H�	NL  *� �K   	� �
�   �� �
�   loc ��K  "G  �
�   (G  �
�   p �NL   �  �
�   8�� �
�   <ctr �
�   @�� �
�   D +K  ^L  =    �~ ��K  �K  �L  =   =    *�� �jL  	`�C     ^L  �L  =   	 *u� ��L  	��e     ^L  �L  =    *i� ��L  	@�e     ^L  �L  =    *%� ��L  	��e     +�� �2  	@�C     /M  /M  =    ^L  +�� M  	 �C     +4� /�   	�'f     ,me 2�   	�'f     +�� 5RK  	�'f     ,wbs 8�M  	�'f     ;  +� :�M  	�'f     O:  ,cnt =�   	�'f     +!� @�   	�'f     -إ C�   +ا E�2  	�'f     +Z� F�2  	�'f     +~� G�2  	�'f     +w� H�   	�'f     +ע I�   	�'f     +� J�   	�'f     +8� M�   	�'f     ,yah UNL  	p'f     +K  �N  =    +�� X�N  	`'f     +� [+K  	X'f     +q� \+K  	P'f     +K  "O  =   	 ,num _O  	 'f     +Ȧ b+K  	�&f     +i� e+K  	�&f     +L� h+K  	�&f     +�� k+K  	�&f     +ܧ n+K  	�&f     +�� o+K  	�&f     +^� p+K  	�&f     +�� q+K  	�&f     +*� t+K  	�&f     ,par u+K  	�&f     +�� v+K  	�&f     +ߢ y+K  	�&f     +{� z+K  	�&f     +9F }+K  	�&f     +\� ~+K  	�&f     +[� +K  	�&f     +K  �P  =    ,p ��P  	`&f     ,bp ��P  	@&f     +>� ��P  	0&f     +K  +U �+K  	(&f     +L� �  	$&f     +ɣ _�   	 &f     �   \Q  =   =    +�� `FQ  	�%f     +� a�2  	�%f     +�� =�2  	�%f     +�� >�   	�%f     +�� ?�   	�%f     +� /�   	�%f     � �Q  �Q  	R  �   �P   .�$ -B     /       ��R  /�  �M  � � 03B     �R  UR  1Uu  28B     �S  3GB     d  3VB     a  3\B     �]   4R� ��R  5� �(�M   .H �xB     ?       �S  3�B     �d  3�B     ja  3�B     �]  3�B     [  3�B     �d   .�� �lB     
       �BS  6vB     �T  1U	�B       7� ��B            ��S  /� �%�   � 
� /�R �5�P  M� G� 8�B     �m  1U�U  .� ��B     r       �1T  2-B     �m  0>B     �T  �S  1U	hB      0MB     �m  T  1U	��C     1T1 8cB     �m  1U	��B     1T1  7%� �hB            ��T  /� �#�   �� �� /�R �3�P  ܀ ր 8vB     �m  1U�U1T1  9&� {B     @      �MZ  /�� /�Q  .� (� :i 	�   �� z� :j �   �� �� +� 
NB  ��:a /M  � ߂ 0�B     �m  DU  1U��1T91Q	��C     1Rv  ;�B     YU  1U�� ;�B     �U  1U	��C     1T	�&f      0B     �m  �U  1U��1T91Q	��C     1Xv  ;B     �U  1U�� ;*B     �U  1U	��C     1T	p'f      ;6B     V  1U	��C     1T	x'f      ;BB     ?V  1U	��C     1T	`'f      0�B     �m  pV  1U��1T91Q	��C     1Xv  ;�B     �V  1U��1T}  0�B     �m  �V  1U��1T91Q	�C     1Rv  ;B     �V  1U��1Tv3$ 'f     " ; B     W  1U	�C     1T	X'f      ;,B     3W  1U	�C     1T	�&f      ;8B     [W  1U	�C     1T	�&f      ;DB     �W  1U	#�C     1T	�&f      ;PB     �W  1U	*�C     1T	�&f      ;\B     �W  1U	1�C     1T	�&f      0fB     �m  �W  1U	9�C      ;�B     X  1U	F�C     1T	�&f      ;�B     BX  1U	M�C     1T	P'f      ;�B     jX  1U	U�C     1T	�&f      ;�B     �X  1U	\�C     1T	�&f      ;�B     �X  1U	d�C     1T	�&f      ;�B     �X  1U	j�C     1T	�&f      ;�B     
Y  1U	r�C     1T	�&f      ;�B     2Y  1U	z�C     1T	�&f      0B     �m  cY  1U��1T91Q	��C     1Rv  ;%B     �Y  1U��1T| `&f     " 0AB     �m  �Y  1U��1T91Q	��C      ;PB     �Y  1U��1T| @&f     " 0uB     �m  Z  1U��1T	TB     1Q9 0�B     �m  .Z  1U��1T91Q	��C      <�B     1U��1T	(&f       .� �~B     |       ��Z  2�B     �m  2�B     �Z  3�B     f  3�B     c  3�B     �_  3�B     �\  3�B     �e   .E� ��B     �       �[  :i ��   � � =�R  ��<  m� k�  .D� ��B           ��\  :lh �	�   �� �� 2�B     ]j  2B     �g  2B     �i  0"B     �m  �[  1U21T2 07B     �f  �[  1U
1T2 0JB     �m  �[  1U21Tv  0\B     �f  �[  1U
1Tv  0oB     �m  \  1U21Ts  0�B     �f  !\  1U
1Ts  0�B     �m  >\  1U@1T� 0�B     �f  \\  1U�1T� 0�B     �m  z\  1U�1T� 6�B     �f  1U
01T�  .d� =OB     �      ��]  2UB     !h  0�B     n  �\  1U01TR 0B     n  �\  1U01T1 0lB     n  ]  1U01T1 0�B     n  4]  1U01TR 0�B     n  P]  1U01T1 0&B     n  l]  1U01T1 0�B     n  �]  1U01T3 3�B     Gf  3�B     �e   .U� 1�B     _       ��]  3OB     Fh   .�� ��B     9      ��_  :i �
�   �� �� :x �
�   N� 4� :y �
�   o� m� =w�  �
�   �� �� 2�B     ]j  2�B     �g  2�B     �i  0B     �m  |^  1T2 0]B     �m  �^  1T2 0�B     �m  �^  1T2 0�B     �m  �^  1T2 0=B     �m  �^  1T}  0dB     �m  �^  1T}  0~B     �f  _  1U| v #@1T~  0�B     �f  ;_  1U| v #�1T~  0�B     �f  __  1U| v #�1T~  8�B     g  1U|�1T~ 1R	�  .�� ]�B            �a  :i `
�   �� �� =d� a
�   7� 5� =�� c�  b� Z� 2�B     !h  0*B     Kd  `  1Ux  0KB     n  `  1U01TR 0uB     n  ;`  1U01T1 0�B     n  W`  1U01T1 0iB     n  s`  1U01T1 0�B     n  �`  1U01TR 0B     n  �`  1U01T1 01B     Kd  �`  1Ux  0`B     n  �`  1U0 0�B     n  �`  1U01T3 3�B     Gf  3�B     �e   .�� A�B     �       �ja  :i D	�    �� 0jB     Kd  \a  1Ux  3�B     Fh   .�� �B     �      �c  :i �
�   � �� >j �
�   :x �
�   �� x� :y �
�   )� � :w �
�   �� �� 25B     ]j  2:B     �g  2?B     �i  0lB     �m  b  1T- 0�B     �m  <b  1U:1Td 0�B     �m  Yb  1U51T2 0�B     �m  qb  1T# 0B     �m  �b  1T}  0;B     �m  �b  1T# 0dB     �m  �b  1T}  0�B     g  �b  1Uv :~ "1T| 1R2 8�B     g  1U}�1T| 1R2  .b� �4B     �      �d  :i �
�   � �� >j �
�   =�� ��  z� x� 2:B     !h  2�B     Kd  0�B     n  �c  1U01TR 0�B     n  �c  1U01T1 2{B     Kd  0�B     n  �c  1U01TR 0�B     n  �c  1U01TO 3�B     Gf  3�B     �e   .>� e�B     t       �Kd  >i h
�   >j i
�   34B     Fh   ?� F�   �B     2       ��d  @# F�   U:i H
�   �� �� =�� I
�   �� �  .� @B            ��d  3�B     �d   .�� �
B     �       ��e  :i 
�   _� U� =r�  
�   ӊ ъ 2�
B     ]j  2�
B     �g  3B     Ri  02B     kh  fe  1Uv1T	`'f      0PB     kh  �e  1U81T	`'f      8mB     kh  1T	p'f       .Ц �
B     6       ��e  2�
B     !h  3�
B     Gf   .r� 
B     #       �f  3�
B     Fh   .-� �i
B            �Gf  2o
B     !h  3}
B     n   Ac� �J
B            �.�) �vB            ��f  B�� �
3xB     S   4ң ��f  Cx ��   Cy ��   Ct ��   >div �
�   >n �
�    4� �g  Cx ��   Cy ��   Cp ��    ?"� t�   �B     �       ��g  Dx u�    � �� Dy v�   w� q� Dn w�   Ӌ Ë /ّ x�   �� }� =͢ {
�   � � :neg |
�   4� 2� =v� }
�   c� a� 0=	B     �m  �g  1U���1T  8j	B     �m  1Us 1T   4� W!h  >i Y�   >a Z/M   4§ $Fh  >i &
�   >a '/M   4*� kh  >i 	
�   >a 
/M   .3� �B     �       �Ri  Dn ��   �� �� Dc ��P  ܍ ؍ :i �
�   � � =Ϸ  �
�   ]� Q� :top �
�   "� � =�T  �
�   ͏ �� =� �
�   C� 9� E�� ��   F�B     n  Di  1U	��C      3�B     �m   .� ��B     n       ��i  :y �	�   B� <� 0�B     �m  �i  1Tv  3B     �m   .]� ��B     �       �%j  :y �	�   �� �� GtB     "       j  ,tmp �B1  ��2�B     �m   82B     �m  1Tv   ?w� �	�  �B            �Wj  Hev �Wj  U '  .�� ��B            ��j  6�B     �m  1U01T0  IFh  �B     �       �k  JTh  J_h  K�B     z       LTh  5� /� L_h  �� �� 2,B     (n  2JB     (n    I!h  qB     �       �`k  J/h  J:h  K�B     �       L/h  �� �� L:h  "�  � 2B     (n    I�g  PB     W       ��k  J
h  Jh  KhB     <       L
h  K� E� Lh  �� �� 2�B     �m    I�f  {	B     /       �zl  M�f  Ŕ �� M�f  A� 7� Mg  �� �� N�f  �  Mg  5� /� M�f  �� �� M�f  � � 0�	B     �m  Ol  1Us 1Tv  6�	B     g  1U�U1T�T1Q�Q1R	�   I�f  �	B     �       �^m  M�f  _� O� M�f  � 
� M�f  Ø �� L�f  w� q� L�f   �� O�f  �   m  M�f  �� � P�f  M�f  G� C� Q�  J�f  J�f  3@
B     �m    0�	B     g  Cm  1Uv 1T} 1R2 8
B     �m  1Uv 1T}   I�R  �B     v       ��m  R�R  US�R   B            M�R  �� ��   T�q  �q  J	T� � 6T��  ��  CT[�  [�  fTj j <T  )'	TL L $ATy�  y�  '9T� � $6T�) �) ?T��  ��  dT� � * 4   ��  S#  �� �*  \B           �� ^�  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  9�  0t  4  e2    �J K   �0  }  ��  (  K B  ڵ  R\  q� �  �� \�  
h0 h   
h1 h  
h2 h  
h3 h  
h4 h  }	 h  
buf 
�  r� 	�   X t    =   ? =�   ��  .N  ^�  2�   }�  7�  �� ;K    	  r�  �   .� $�  O� )�   �  �  �        �  �   �  1   �  �  K   R   1    �  ��  ,N  �  t  oS  	'�  dS  (	)O  � 	+
O   � 	,�  @�  	-
�   >z 	.
�   �  	/R   �H  	3_    �   _  =    �  	�� 	7_  	�� 	8K   �� �  	 (f     �  �� �   	�'f     � D\B           �s  j� D�  �� �� �� F�  ��~i GK   � � s  �B      0  R	<  �  4� 2� �  i� W� 0  �  ��~�  �B      �B     L       ?$�  �  5� 3� �B     L       �  ^� X� �  �B     �  T|    �B     �  �  U��~Ts Q9 �B       �  U��~T��~ B         U��~ +B       %  U��~ 8B       U��~   ~B       U  U��~ LB     +  U��~T��~   �� 9�  !�� 9-�  !�O  9G_  "buf ;
�   �  �   �  =    #ͨ �   �  !t &�  "i !	�   $��  "	�    %�� �� 
B%  '	%�� �� %%M� M� $%� � !%-� -� # �   ��  S#  � �*  ^B     '       
� ��  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  ڵ  RI  	�  �   	q  y  �   =� �  ��  .�  ^�  2M   }�  7S  �� ;K    
	�  r�     .� $  O� );         �      �          1   ;     K   R   1      ��  ,�  A  U  	� A  M  u  =     ۨ (e  %� Z1   B            �  wad Z   �� �� 82  Z-K   � � �< [R   %� !� � [$1   b� ^� �B     U�UT�TQ�QR�R  �� UyB            �^  wad U   �� �� B     U�U  � 5   ^B            ��  �> 5�   �� ؝ ��  7    i 8	�    lB     �  �  U	��C      yB     U�U  � � ! %   4�  S#  ,� �*  �B     k       %�  �  �)  �=   ,	  0t  P   e2    �  �0  }  int ^&  ��  D   ^   J�   D   �C  
D  ���� �C  N�   ڵ  R�   �   1  	�  s   	q  �   �   
�1  @y  Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2s   8;:  5s   < �K 8"�   	�  K�  y  	�  L�  	�  M�  =� �  ��  .�  ^�  2}   }�  7�  �� ;^    	!  r�  6   .� $G  O� )k   0  0  �    �  !  G  0   <  1   k  0  ^   �   1    M  ��  ,�  q  �   oS  	'�  dS  (	)�  � 	+
�   � 	,0  @�  	-
s   >z 	.
s   �  	/�   �H  	3    �     =    �  	�� 	7  	�� 	8^   �
 	�   �B     k       ��  �   �   C� ?� p !	s   � {� �B     !       �  ��  ��   �� �� �B     �  �B       �  U	WB     T|  �B       U|   �B       U	��C     T1  ��  ��  
+��  ��  d� � 	:��  ��  % P   ��  S#  ͩ �*  �B            �� ��  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  �   	int �K 8"T   
�  K  �   
�  L  
�  M  9�  0t  9  e2    �0  }  ��  -  K   J�  D   �C  
D  ���� �C  Na  ڵ  RU  K   �  7�  � �   }  <�  ;�  1^  o�  f~  ��  	 ��  (�  K   /!  ��   [r  �4 #�  �   �  
��  ��   
�\  ��  
�  �K  �  
��  ��   
��  ��   
2�  ��  
��  ��   
Ɇ  �!  
��  ��   
��  ��   
�h  ��   
rK  ��   
l�  ��   
]�  ��   
��  ��   K   	"'  ��  WH  �~  �O  �m  ��   �  ��  ��  	 =� 
3  ��  
.h  ^�  
2�   }�  
7!  �� 
;K    
	�  r� 
 �   .� 
$�  O� 
)�   �  �  �    '  �  �  �   �  1   �  �  K   R   1    �  ��  
,h  �  oS  '  dS  ()c  � +
c   � ,�  @�  -
�   >z .
�   �  /R   �H  3s    �   s  =    �  
�� 7s  
�� 8K   '	�  �� *�   �� +�   2� ,�    �   �  =    � -�  0	  � 2�    >z 3�   � 4c   �� 5�  y  =	 �i     �  >	(f     ĩ BU  	(f     s  ?�  4h  A�   � B�    [  �  �  =    �  թ C�  	`�C     � Jn#B     �       ��  4h  J'�  
� � i L	�   X� V� C� M	�   ~� |� �#B     �  2  Us h�C     " �#B     b  J  Uv  �#B     b  b  U|  �#B     n    Uv T4 �#B     z  U	��C     Q	��C     R} X	��C     Y�H  Z �"B     �       �Z  i K   �� ��  ;#B     +       3  ȩ .K   ޟ ܟ Q#B     �  Us   !�"B     �  #B     �  T1Qv   �q  ��"B            ��  � ��   
� � �"B     :  �  U�U "�"B     �   } ��"B     K       �K  C� ��   I� C� �O  �s  �� �� �"B     z  #  U	��C     Ts  #�"B     �  T8Q	��C     R
�  $��  �R   o"B            ��  � ��   +� '� %tag �'�   h� d� |"B     :  �  U�U #�"B     �  T�l�  $� ~R   �!B     �       ��	  C� ~�   �� �� %tag ~'�   � � ��  �!  `� X� �O  �s  �� �� �!B     z  d	  U	n�C     T}  9"B     �  �	  Uv T| Q	��C     R
� C"B     �
  �	  U}  Q"B     �  �	  T| Qs `"B     �	  U}   { Vn!B     f       ��
  �O  VK   � � `5 V*R   N� H� c X	�   �� �� l Ys  ֣ ԣ &~� l�   c
  ' �!B     z  �
  U	)�C     Tv  !�!B     �  �!B     �  �
  Q|  �!B     z  �
  U	D�C     Rv  "�!B     �   $�} E�   E!B     )       �:  �O  E K   �� �� ^!B     z  U	�C     Ts   $�{ 2�   !B     &       ��  � 2�   Q� K� i 4	�   �� �� *!B     �  �  Uv  ?!B     z  U	��C     Tv   (j  �     )�  �   *+� s  +i 	�   ,*ȩ 	�     - � ��   � B            �.� ��  &B     \      ��  /��  ��   � � n� ��  ��0+� �s  .� &� 1i �K   �� �� 0� ��  � ݥ 0�� �	�   X� V� 0� �	�   }� {� 0u� ��  �� �� 0�� ��  � � 0�� �	�   �� �� 2�  FB     p  ��  3�  ا ֧ 4p  5�  �� �� 5�  ;� 5� 6�  �B     .       t  5�  �� ��  KB     �  �  Uv  $ &T( _B     z  �  U	��C      �B     �  �  Tw # !�B     �    <B     �  �  Us  SB     �    U	��C     Ts  {B       =  T	/PB      �B     �  ^  U@T1Q0 �B       |  Us T| �B     �  �  U} T0Q��R< �B     #  �  U��T	��C     Q4 �B     #  �  U��T	��C     Q4 	B     z     U	��C     Ts  B     �  B  Us T1Q0 3B     �  l  U} Q| Rs  $ & J B     /  �  UsXTpQ8 T B     �  �  U|  !e B     �     7	� W�  8�� W �   9�� Ys  :i ZK   ,9?� s�     .� FK   �B     6       �a  ;s F)a  �� �� 0��  KK   � � 1i LK   [� W� !B     ;   �   <�  � B     �       �b  3�  �� �� 5�  � � =�   � B     C       �  5�  L� H� � B     �  �  U|  � B     G  Us T| Q8  >�  � B     0       3�  �� �� ?� B     0       =�  5�  ê �� !B     G  Uv(T| Q8    @� � _@��  ��  0@��  ��  7@� � 	7	@� � 	6@�� �� 	<	@�� �� p@%� %� 
KA~� ~� l@� � ?@K� K� 	=	@m�  m�  @@� � 
A@��  ��  d@:�  :�  @�^ �^ #@-` -` @�` �` @� � @� �  �	   ��  S#  �� �*  �#B     /      }� ~�  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  
K   	"f  ��  WH  �~  �O  �m  ��   �  ��  ��  	 0t  r  e2    �0  }  ��  f  ڵ  R�  ٪ ('  >z )�    m� *  tag +�   id ,�   �H  -  s�  .    R   �  � /�  82	J  >z 5
�    �� 8  �� :J  0   Ī <  X� @r  	(�i     P  r� �K   )B     
       ��� ��   �(B     ,       ��  �� �J  � � m�  ��   � �  K� ��(B     *       �_  ptr �R   N� F� m� �%  �� �� �� �J  � �� �(B     �	  U	��C       �� �i(B     V       �:  ptr �R   z� t� tag �"�   ̬ Ƭ � �-�   � � ��  �7�   q� k� �� �J  í �� �(B     �	    U	$�C     T| Q}  �(B     �	  U	P�C     T| Q}   [ ��'B     q       ��  �� �J  � � /(B     �	  �  U	��C      E(B     �	  �  U	��C      a(B     �	  U	��C       �� oF'B     �       ��  f o  A� ;� �� qJ  �� �� d'B     �	  4  Uv T	%�C      �'B     �	  _  Uv T	W�C     Qs  �'B     �	  �  U	�C     Tv  �'B     �	  �  U	7�C     Tv  �'B     �	  U	h�C     Tv   Ϊ H�&B     �       ��  }� I�   �� �� �� J�   
� � �� LJ  X� V� �&B     �	  H  U	%�C      �&B     �	  s  U	B�C     Tv Q|  �&B     �	  �  U	W�C     Ts  'B     �	  �  U	��C      !'B     �	  �  U	��C      ;'B     �	  U	��C       E} *4&B     P       �s  }� +�   �� {� �� ,�   ӯ ͯ �� .J  %� � �H  /J  r� p� z&B     �   � �R   &%B           ��  >z ��   �� �� tag ��   #� � m� �
R   s� m�  P �
�   ñ �� ' �J  �� �� �� �J  !� � �� �J  F� D� �1  �J  s� i� ��  �R   � � s%B     �	  n  U	��C     T|  �%B     �  �  Uv( �%B     �	  U	��C       � ~{$B     �       �	  ptr ~R   � 	� �� �J  v� r� �  �J  �� �� �$B     �	  U	��C       � a'$B     T       �n	  �� cJ  � � >z d
�   �l5$B     �	  U�l  a� G�#B     7       ��	  \� Gr  U�� IJ  %� !�   ��  ��  7 F�  F�  b!�E �E   ��  ��  d!      �C �C #     ��  S#  ]� �*  )B     �       �  ��  �)  �=   ,	  ^&  �  �1  @�   Q  �    �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2�   8;:  5�   < �   1  int �K 8"T   	�  K  �   	�  L  	�  M  0t  -  e2    �0  }  ��  !  ڵ  RI  =� m  ��  .�  ^�  2/   }�  75  �� ;K    
	�  r�  �   .� $�  O� )   �  �  �    a  �  �  �   �  1     �  K   R   1    �  ��  ,�  #  U  K   "�  ��  WH  �~  �O  �m  ��   �  ��  ��  	 
 	�  wad a   }_    8� �  	� #  �  Y	��e     H� E1   )B     2       ��  wad E �  b� \� 82  E2K   �� �� �< FR   � � � F)1   Z� R� T� H�  �� �� ��  I1   9)B     �  �  T	�T����Q0 Q)B     �  U�QT1Q�R  �  '� 8Q)B            �  wad 8*�  � � T� :�  z� r� ^)B     �  g)B     �  U�U  k� !�  g)B     P       ��  �> !*�   ݶ ٶ ��  #�  � � }_ $  T� P� t)B     �  �  U�UT	P�B      �)B       �  U T1Q0 �)B       Uv   VL VL ��K �K �5L 5L Y� � 7	�/ �/ [� � 6�] �] 	! m	   ��  S#  �� �*  �)B     �        ��  �)  �=   ,	  int ^&  9�  �� �  }  �  e2  �1  @  Q     �   	1   62  #	1     &	1   �5  )	1    �@  ,	1   (.  -	1   0*  2D   8;:  5D   <   1  	  �K 8"~   
�  K+    
�  L+  
�  M+  0t  w     �J p   �0  ��  I  K \  p   J�  D   �C  
D  ���� �C  N�  ڵ  Ro  	�  p   !�  �p   �  ��  S�  ��   �F  '�  *	L  *� ,�   "G  C	D   (G  CD   �]  CD   :G  CD    �U  D   (	�  ��  ,	D      -	D   &: 4�  �9 9�  �= Y�   �  �   �  �  �  �  D   D   D   D    �  ]< ZX  
��  �  
�\  ��  
�  �b   
��  �D   
��  �D   
2�  ��  
��  �D   
Ɇ  ��  
��  �D   
��  �D   
�h  �D   
rK  �D   
l�  �D   
]�  �D   
��  �D   
: 	�  
O: 	�  
k: 	 �  
�: 	!�  
]: 	"�  
K; 	&�  
�; 	'�  
�; 	(�  
�; 	)�  
< 	*�  
�: 	.�  
; 	/�  
<; 	0�  
r; 	1�  
�; 	2�  
�  
D   
q  
j    
��  %  t�   D   	|  �  �  =   �' 	�  
��  1�  
]  4�  �  �  �  =   � 	�  
Zy  8�  �  �  =   =   � 	�  
��  ;�  Ʃ  Qp   	
    ,  =     	  
�  W,  D   M  =    
N�  %=  
��  '�  =� q  ��  .�  ^�  23   }�  7�  �� ;p    	�  r�  �   .� $�  O� )!   �  �     e  �  �  �   �  1   !  �  p   K   1      ��  ,�  '  oS  'E  dS  ()�  � +
�   � ,�  @�  -
D   >z .
D   �  /K   �H  3�      �  =    9  
�� 7�  
�� 8p   
UK 
�  {    ,	ȓe     �� 0D   	(f         =    		  1� 3  � 1234567890-=	qwertyuiop[]�asdfghjkl;'`�\zxcvbnm,./�*��������������                                 � �� �                  �� �  	��C     �� Rf*B            �Ѱ �)B     �       ��  u L  �\ǭ 	D   �Xkey w   �W�  �)B      �   	s  	  �� �� �  �� �� �  	  ٷ շ   	  *B        *�  -	  � �   �)B     X	  �  !U�X!T�W  8*B     d	  �  !U�\ "a*B     d	  !U�\  #u� 	  $ǭ #D   %key :w   &�q 		D    '� �w   :	  (key �1w    '�� �w   X	  (key �1w    )�� �� )i�  i�  � �   ��  S#  ʳ �*  g*B     �      �	 4�  T   A   F   - 1   ,	  1  M   e� A   �� �)  �F   0t  �   e2  ޱ �     �J �   �  �0  }  int ^&  ��  u   H� �   K �   	�   J  
D   
�C  
D  ���� �C  N�   ڵ  R�     �   ?  F    N�  %/  ��  'W    �  �   q  u  {  M   �1  @  Q  {   �   	i   62  #	i     &	i   �5  )	i    �@  ,	i   (.  -	i   0*  2�   8;:  5�   < �K 8"�  �  K    �  L  �  M  	�   	;�  
�  
� 
| 
7	 
 
�
 
` 
� 
� 
� 	 � 	F:  � 
.�  I� \�  �    ��  �{  �\  �  �  ��  �  ��  ��   ��  ��   2�  �  ��  ��   Ɇ  �W  ��  ��   ��  ��   �h  ��   rK  ��   l�  ��   ]�  ��   ��  ��   	�   "�  
��  
WH  
�~  
�O  
�m  
��  
 �  
��  
��  	 t�   �   �  �  �  F   �' �  ��  1�  ]  4�  �  �  
  F   � �  Zy  8
  *  1  F   F   �   ��  ;1  Ʃ  Q�   B  N  d  F     S  �  Wd  UK 
�  �   9�  n� 4�  82  6�    �� 7�    `� 4:9  J� <�    z� =�   �� >�   �� ?�   �� A�   red D�  �� E�  �� F�  $^� G�  , �� J�  	@,f     �� K�   	ԓe     1� L�   	8(f     g  N�  b O�    g P�    r Q�    a R�      {  �  F   � ��  U�  	@(f       [	0(f     !� \W  	((f     �  `		$(f     �  e		0�i     �  p	Гe     �  q	̓e       u	 (f     w	�  r y   g z  b {   Q� |i  �   �  F   � 9� ��  � �# ��.B            ��  4� �   U � �� � ��.B            �5  ڈ �3�  U  �� ��.B            ��  �4 �{  �� �� �.B     i  U�U  ~� ��� � T� \�   �.B     I       �r  !r \�   ׸ Ѹ !g \#�   '� #� !b \*�   d� `� "< ^	�   �� �� "�< ^�   ޹ ع #�< ^�   $i _	�   0� ,� "g  `�  m� g� %�.B     u  U	��C       � >>.B     ]       ��  @� >W  պ Ϻ $i @�   (�  �   1/.B            ��  !scr 1W  �� ��    Y-B     �       ��	  $y 	�   ƻ Ļ "�� 	�   � � "W� �   � � "<� �   a� ]� "d� �	  �� �� "�� �	  �� �� &�-B     H       �	  $i �   � � %�-B     �  Uv Tt Qq   '/.B     �   �   (�
 �)� �S-B            �
  'X-B     �   (� �)l� �8-B            �\
  *E-B     �  'R-B     �   )} ��+B     �      ��  +i �	�   6� 2� ,�� ��   -#,B     �  �
  U	`�C     T
�Q
�R
�X
�Y  -e,B     �  �
  U	��C      -,B     �  $  U	!�C     T
@Q� -�,B     �  H  U	S�C     T1 *�,B     �  *�,B     �  -�,B     �  �  U
 �T1Q0 *!-B     �  '8-B     �   )� ��*B     �       ��  .out ��  z� l� .in �*�  (�  � /Z� �2�   Q+i �	�   �� �� +j ��   � �� +k ��   Q� M� +c �{  �� �� +pix ��   � � +r ��   J� F� +g ��   �� �� +b ��   (� &�  �   )�� �g*B     a       �L  .out � L  r� l� .in �/�  �� �� /Z� �7�   Q+i �	�   6� 0� +j ��   �� �� +c �{  �� �� +r ��   �� �� +g ��   �� �� +b ��   K� G�  �   05  �.B            �1� � 2     1� � 1Ѱ Ѱ W1� � 7	1m�  m�  @1��  ��  d1��  ��  %1� � (1� � 61��  ��  A1�� �� �    �  S#  ܳ �*  �.B            � 3�  e2    �J K   �  ,	  �0  }  int ^&  K ?   UK 
�   u   �   	x,f     �  �.B            �   	��      �   
R    �.B       �   U�<$ /B        ��  ��   Գ Գ  �   �  %� ˹ �*  p          � ��  �)  �9   ,	  ^&  �  �1  @�   Q  �    �   	-   62  #	-     &	-   �5  )	-    �@  ,	-   (.  -	-   0*  2�   8;:  5�   < �   1  �   	int �K 8"P   
�  K  �   
�  L  
�  M  0t  .  e2  ޱ A    �J G   � 9   �0  }  ��  "  H� 5  K H  j� T  �� N   � (  x �    y 	�   ��  �     �   �9 �   � 
n  �< 	  �� 

n    n  `� �  �� 	R  x 		�    y 	�    q� 		.  K� 	�  r 	n   g 	n  b 	n  a 	n   �� 	^  9�  �� �� std  �  &� AA�  
A  
�u  
��  
��  
��  
�  
�!  
�7  
��  
��  
��  
��  
��  
�  
�;  
�\  
�n  
�z  
��  
��  
��  
��  
�  
�)  
��  
��  
�D  
�_  
��  
�u  
��  
��  abs f-� ?	  �  ?	   abs T�� N	    N	   abs NE� �  "  �   abs J�� �  <  �   abs F#� �  V  �   abs =�� �  p  �   abs 8W� @   �  @    div 
�.� u  @   @     �   &� AA�  
��  
�D  
�_  
�u  
��  
��  
��  div 
�#� �  �  �    P� A  9� �    rem �    Q�   Z� u  9� @    rem @    [� M  ; �  9� �   rem �   ξ �  �� I�   �  �   �  Z� J�   �  �   �M '�  �     �� �   � (�   !     �� )@   7     �� VN   a  a  a  -   -   h   g  n  �   �  a  a   div aA  �  �   �    � M�   �     � bu  �  @   @    �� g�   �    -    N� m-   	  	    -      &�    �� h�   ;  	    -    �� X\  N   -   -   h   ]� N#n  �    � 5�   � 7�  G    �� +�  �    �   �   � .@   �    �  �    �� 09   �    �  �    C O�        l� n-   #  �   #  -      �� i�   D  �      � c	�  _  �  �   �� *�  u      � /�  �    �  �    _� 1�  �    �  �    2� �� ,�  �    �   �  � -�  �    �   '�  +�  .\  3A  4u  abs ]�   7	  �    6!	  �� 6�  G� 6�  6  6"  6<  6V  6p  7�  8  9!  :7  <�  <�  <�  >�  @�  C�  D�  E  G;  Hn  Jz  K�  L�  M�  N�  P  Q)  R� "  �� �  {� I� \
  b
   �   �� �� w
  �
   �   �    �� !�� �
  �
   �   	� *�� �
  �
   �     c� ;�� �
  �
   �     !�� L5�   �
     �  G    !�� P\�     %   �  G    � Z?� :  J   �  G      !�� d9� �   c  i   �   !n� h��   �  �   �  G    !:� }O�   �  �   �   !u� �D�   �  �   �   "g� �   "� �  #num �G   $T    :
  	  %�� %4�   � %  +  &6  4
   |� �  x z   y z  ��  z    z  �  �  �4 �  e� �  lt �  t'� u� �       (�   �  )9   _ � 6  �� � g  �� !:
   t #�  y� $�   U &-�  �G� ("  �׺ )  ��� *  ��� ,�   ��� -R  ��� /  � (� �  0� �   � �  msg �  "8 �  (G  �    � g  (A  �  )9    *�� �  	 -f     *7� G   	-f     *�� G   	-f     +L� 	*  	 -f     �  +� �  	�,f     
UK 
R  �  ,=� @            ��  -�  @     @            �.�  �� �� .�  �� �� -  @     @            /,  
�,f     �   0��   1"� ��   1�� ��    2� ��0B     $       �d  3�4 �%  �� �� 4
1B     M  V  5Us,5T�U 61B     Y   7�� ��   �0B     2       ��  8ǭ ��  U8�� �,�  T9�0B     !       :E� �A  M� K�   �   .  7}K y
�  �0B     &       �  *�� {�  �`;ms |�  �h 2JK t�0B            �G  <ms t�  t� p�  2� ^�/B     �       ��  ;msg `�  �H40B     e  �  5U�H =<0B     K  =J0B     q  4Q0B     }  �  5U0 4p0B     �  �  5Q�<$ =|0B     �   2Գ R�/B     E       �K  4�/B     M  /  5U	�,f     5T	��C      >�/B     �  5U	�,f       ?L� G/B     �       ��  3ǭ G�   �� �� 3�� G5G   !� �� @key I.  |� z� :E� KA  �� �� A�  /B     @  I&.  �� �� >a/B     �  5U�T   B�  .    Ckey  4G    �    D�  ,  6  EY    F  V� G  M  G,   H�� �� H� e� <H� Y� 
HS� � 9Hc� c� K#H�� �� Hm� E� 6H� �� 8	H/� /�  �   Z�  � ?� � 1B     u       � e2    �  � N   ,	  �0  }  int ^&  N� �N   j� B   �� 4q   (� �   0� }    � }   msg }   "8 }   (G  }     � �   (� 
�� F1B     D       �\  	pid 
}   �@	msg 
.�   � 
m }   �`"8 }   �X(G  }   �P Y� 
� }   1B     1       ��  	msg (�  �P4� }   �` �    �   <�  � �� � �1B     E      � 0t  9   e2  ޱ L     �J _   �  � r   ,	  �0  }  int ^&  ��  -   H� @   K S   j� f   � (7  x �    y 	�   ��  �     �   �9 �   � 
�   �< 	7  �� 

�     �   `� �   @� �  ��  �      �   bpp 	�   �9 �   
 �� I  �� �  x 	�    y �    q� 	�  D� �  pos �   >z �   � �  K� 5  r �    g �   b �   a �    �� �  	'�� �  �� (�   >z )�   $� *�   82  +�   
 
�  �  r    1  �  �� ,A  �)  �r   std  r  &� 
A
A�    �C  ��  ��  ��  ��  ��  �  �W  �r  ��  ��  ��  ��  �  �7  �I  �U  �g  ��  ��  ��  ��  �  �~  ��  �  �:  ��  �P  �p  ��  abs 	NE� �  �  �   abs 	J�� �    �   abs 	F#� �  "  �   abs 	=�� w  <  w   abs 	8W� �   V  �    div �.� C  �   �     � 
�  &� 
A
A  �~  �  �:  �P  �p  ��  ��  div �#� ~  w  w    	P�   9� �    rem �    Q� �  	Z� C  9� �    rem �    [�   	; w  9� w   rem w   9�  ξ O  �� I�   �  �   �  Z� J�   �  �   �M '�  �  �   �� �  � (�   �  �   �� )�     �   �� V�  6  6  6  �  �  =   <  C  �   W  6  6   div a  r  �   �    � M�  �  �   �  � bC  �  �   �    �� g�   �  �  �   N� m�  �  �  �  �   �  &�  �  �� h�     �  �  �   �� X7  �  �  �  =   ]� N#I  �    � 5�   � 7g  _    �� +�  �  �  �   �  � .�   �  �  �  �    �� 0r   �  �  �  �    C O�   �  �   l� n�  �  �  �  �   �  �� i�     �  �   � c	~  :  w  w   �� *w  P  �    � /w  p  �  �  �    _� 1�  �  �  �  �    2� �� ,�  �  �  �   �  � -�  �  �  �   �� '�  +�  .7  3  4C  abs ]�   	  �    6	  6�  6�  6  6"  6<  7�  8�  9�  :  <�  <W  <V  >r  @�  C�  D�  E�  G  HI  JU  Kg  L�  M�  N�  P�  Q  �� �b� �=B            ��
  `5 �'�
  �H src �8�
  �@82  �H�  ��!�� ��
  �`!�� ��
  �X"�=B     �       #i �
�   �l">B     �       #j ��   �h   =  �   $� � � p<B     ?      �V  `5 ��
  �X src �-�
  �P82  �=�  �H
� �L�  ��!�� �	�   �h!�� �	�   �d!�� �	�   �`"=B     �       #i �
�   �l  $� �n� �;B     �       ��  `5 ��
  �X src �-�
  �P82  �=�  �H"�;B     �       #i �
�   �l"�;B     �       !�� ��   �h   $�� �e� 
:B     �      ��   x ��   �\ y �&�   �X��  �-�   �T  �8�   �P c1 �N5  �L c2 �`5  �HG� �o�
  � "q:B     #      #j ��   �l  $�� �Q� �9B     W       ��  � �"�  �` c1 �65  �\ c2 �H5  �XG� �W�
  �P $�� �� I8B     j      ��   x ��   �\ y ��   �X��  �%�   �T  �0�   �P c1 �F5  �L c2 �X5  �HG� �g�
  � "�8B     %      #j ��   �l  $^� ��� �5B     J      ��   x ��   �� y �!�   �� w �(�   �� h �/�   ��"8 �;7  ��G� �L�
  ��!� ��  �B!�� �
�   �_!�� ��   �X!F� ��   �l!�� ��   �h!�� ��   �T"�6B     �      #i ��   �d"�6B     ~      #j ��   �`"�6B     K      !82  ��   �P    $�� ��� �5B     Q       �:   x ��   �l y ��   �h��  �!�   �d  �,�   �`�� �B5  �\G� �U�
  �P $�� ��� �4B           �;   x ��   �L y ��   �H��  �!�   �D  �,�   �@ r �<�   �� g �G�   �� b �R�   ��G� �`�
  �!I� ��   �h!�< ��
  �`"5B     �       #i ��   �l"65B     l       !� ��   �\!��  ��   �X   $�� ��� M4B     I       ��  � ��  �`�� �*5  �\G� �=�
  �P %�v ��� �   4B     .       ��   num ��  �X#x ��   �l %� ~��   �3B     [       �  � ~�  �PN}  ~*�  �H R� &�� p � �
  O3B     u       �n  �� p/�  � �� p=�  �X!G� q�
  �h $�� ]�� j2B     �       ��  `5 ]�  �X src ])�  �Pr� ]5�  �H!� c	�  �h!�� d	�  �` $R� I�� �1B     �       �H  `5 I�  �X c I.�   �Pr� I8�  �H!� R	�  �h!�� S	�  �` '�� 5G� �1B     8       �`5 5�  �h c 5.�   �dr� 58�  �X  �   ��  � �� �            �' 0t  5   e2  ޱ H     �J [   �  � n   ,	  �0  }  int �   ^&  N� �n   ��  )   H� <   K O   j� b   �� 4�   �� �   � (^  x �    y 	�   	��  �   	  �   	�9 �   	� 
�   	�< 	^  	�� 

�     
�   `� �   �� �  x 	�    y �    q� 	p  D� �  pos �   	>z �   � �  K�   r �    g �   b �   a �    �� �  1    �)  	�n   9�  �� �� std     &� AAP  
�  
��  
�  
�,  
�B  
�e  
�{  
��  
��  
��  
�  
�.  
�I  
�{  
��  
��  
��  
��  
��  
�  
�-  
�M  
�c  
��  
�  
�W  
��  
��  
�  
��  
��  
�>  abs NE� 9  |  9   abs J�� 7  �  7   abs F#� X  �  X   abs =�� 2  �  2   abs 8W� �   �  �    div 
�.� �  �   �     � s  &� AA  
�  
��  
��  
��  
��  
�  
�>  div 
�#�   2  2    P� �  	9� �    rem �    Q� s  Z� �  	9� �    rem �    [� �  ;   	9� 2   rem 2   ξ �  �� I�   %  %   
+  Z� J�   B  %   �M 'X  X  _   �� 
!  � (�   {  _   �� )�   �  _   �� V�   �  �  �  &  &  �   
�  
�  �   �  �  �   div a�  �  �   �    � M    _   
  � b�  .  �   �    �� g�   I  _  &   N� m&  i  i  _  &   
o  &�  o  �� h�   �  i  _  &   �� X�  �   &  &  �   ]� N#�  �    � 5�   � 7�  [    �� +X    _     
  � .�   -  _    �    �� 0n   M  _    �    C O�   c  _   l� n&  �    �  &   
v  �� i�   �    o   � c	  �  2  2   �� *2  �  _    � /2  �  _    �    _� 1    _    �    2� �� ,7  7  _     �  � -9  Y  _     '  +,  .�  3�  4�  abs ]�   �  �    6�  6b  6|  6�  6�  6�  7B  8e  9{  :�  <W  <�  <�  >�  @  C.  DI  E{  G�  H�  J�  K�  L  M-  NM  Pc  Q�  R� 
d  �� ?  {� I� �	  �	  ?   �� �� �	  �	  ?  �    �� !�� �	  �	  ?   	� *�� �	  �	  ?  J   c� ;�� 
  
  ?  J    �� L5� J  8
  C
  ?  [     �� P\� J  \
  g
  ?  [    � Z?� |
  �
  ?  [   J    �� d9� �   �
  �
  ?    n� h�� J  �
  �
  ?  [     :� }O� J  �
  �
  ?    u� �D� J      ?   !g� ��   !� ��  "num �[   #T J   
|	  ?  
P  $�� 4� �  !�H  	�   !s�  
�  "obj J  %�� G� �  �  �   #T J   
U  �  � �  
�  &�  v	   |� Y  x �    y �   	��  �   	  �   	�  �   	�4 Y  	e� �   l	t �   t'� u� R  �    (  i  )n   _ � �  �� � 4  	�� !|	   	t #�   	y� $i   	U &-  �	G� (d  �	׺ )^  �	�� *^  �	�� ,�   �	�� -�  �	�� /�  �*�� ��        �    '�� b� -      +�
  S  �GB     -      ��  ,Y E  �H-pos h[   �D.�� n�  �h/obj rJ  �X0�GB     	       �  .v� jJ  �P 1�GB     8       /i p[   �d  +�	  �  �FB     �       �  ,Y E  �H-obj *J  �@.=� +�  �X 2�  ,  6  3Y �   4  �� Y  �FB     "       �b  5,  �h +
  �  �FB     "       ��  ,Y E  �h-pos L[   �d 6C
  �   FB     �       �  ,Y E  �X-pos P[   �T.�� S�  �h1FFB     8       /i U[   �d  6�
  %  �EB            �2  ,Y E  �h 7�	  @  S  3Y E  3m� �    82  c� v  �EB     -       �  5@  �h 7�	  �  �  3Y E   4  !� �  �EB     -       ��  5�  �h 9�� ~*� �DB     &       �  :\� ~J  �h-win ~(  �` 
u    9�� p� �CB     �       ��  -win p"  �H:�� p2�  �@;�  /i u�   �l1-DB     c       .�� v
�  �P   <_� g	�� J  /CB            ��  -win g  �h:�� g/�  �` 9� \w� �BB     �       �>  -win \  �H:�� \.�  �@;�  /i ]
�   �l1�BB     p       .�� ^
�  �P   9�� MG� �AB     �       ��  -win M  �X1�AB     M       /i Q
�   �l  9E� Cm� +AB     �       ��  -win C   �h =e� ?� �@B     6       ��  -win ?  �` 9� :S� �@B     C       �%  -win :  �X 2   6  I  3Y 
  3m� �    8%  8� l  vEB            �u  56  �h <�� %	�   �?B           ��  :y� %"�  ��/win '
  �X.t )�   �P.G� -d  �� 
i  �  2    �     3Y 
   8�  �� #  �DB     �       �,  5�  �h 2E  =  G  3Y �   4,  V� j  �DB     2       �s  5=  �h =�� !H� �?B     0       ��  :L� !�   �`:�< !(�   �\ =� �� Q?B     /       ��  :L� �   �` >�� 
q� �   ?B     D       �G  :@� $�  �P:׺ 4G  �H:�� JG  �@/h �   �` 
�   ?�� 
z� �   �>B     >       �:@� $�  �P/h �   �`  Q    ��  �HB     �IB     �. ../src/gfx/sse2.asm NASM 2.13.02 ��HB              �   ��  �  � � �IB     �       8/ ^&  �)  �@   ,	  9�  �� �� std    &� AAe   �  ��  �-  �J  �`  ��  ��  ��  �  �!  �=  �X  �s  ��  ��  ��  ��  �  �  �>  �^  �~  ��  ��  �!  �l  ��  ��  �M  �  �&  �o  	abs NE� N   �  
N    	abs J�� h  �  
h   	abs F#� v  �  
v   	abs =�� G   �  
G    	abs 8W� -   �  
-    div �.� �  
-   
-     � �  &� AA"  �!  ��  ��  �  �&  �M  �o  div �#� !  
G   
G     P� �  9� �   rem �   int Q� �  Z� �  9� -    rem -    [� �  ; !  9� G    rem G    ξ �  �� I�  C  
C   I  Z� J�  `  
C   �M 'v  v  
}   �� �  1  �  � (�  �  
}   �� )-   �  
}   �� V�  �  
�  
�  
4   
4   
�   �  �  �    
�  
�   div a�  !  
�  
�   � M7  7  
}   �  � b�  X  
-   
-    �� g�  s  
}  
4    N� m4   �  
�  
}  
4    �  &�  �  �� h�  �  
�  
}  
4    �� X�  
�  
4   
4   
�   ]� N#�  
�   � 5�  � 7  
   �  �� +v  8  
}  
8   7  � .-   ^  
}  
8  
�   �� 0@   ~  
}  
8  
�   C O�  �  
}   l� n4   �  
7  
�  
4    �  �� i�  �  
7  
�   � c	!  �  
G   
G    �� *G     
}    � /G   &  
}  
8  
�   _� 1F  F  
}  
8  
�   2� �� ,h  h  
}  
8   �  � -N   �  
}  
8   '-  +J  .�  3�  4�  abs ]�  �  
�   6�  6w  6�  6�  6�  6�  7`  8�  9�  :�  <l  <  <�  >!  @=  CX  Ds  E�  G�  H�  J  K  L>  M^  N~  P�  Q�  �� )�� ;JB            ��  p )�  �h@   �` �� #��  JB            �  p #�  �h �� �� JB            �@  p �  �h@   �` �� �� �IB            �p  p �  �h �� �� �  �IB     )       ��   >z (@   �h !�� �� �  �IB     )       � >z &@   �h  %U�B   :;9I  $ >  :;9   :;9I8   I  $ >  4 :;9I?<  	.?:;9'I@�B  
 :;9I�B  �� 1  ��1  �� �B  . ?<n:;9  . ?<n:;   %�B  $ >  $ >  >I:;9  (   (    :;9I  4 :;9I?  	. ?:;9'@�B   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  (   :;9  I  ! I/  ! I/       '   I  :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  ":;9  # :;9I8  $ :;9I8  %:;9  &:;9  ' :;9I8  ( '  )(   *'I  +4 :;9I?  ,4 :;9I  -4 :;9I  .4 G:;9  /4 :;9I  04 :;9I  14 :;9I  24 G:;9  3.?:;9'@�B  4��1  5�� �B  6�� 1  7�� �B1  8 :;9I  94 :;9I�B  :��1  ; :;9I�B  <.?:;9'   =4 :;9I  >4 :;9I  ? :;9I�B  @ :;9I  A4 :;9I�B  B���B1  C.?:;9'I@�B  D. ?:;9'@�B  E.1@�B  F4 1  G4 1�B  H  I. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  (   :;9   :;9I8       I  ! I/  ! I/  '   I  :;9   :;9I   :;9I  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  " <  #:;9  $ :;9I8  %4 G:;9   %�B  I  !    I  $ >  4 :;9I?<  4 G:;9   %�B  $ >  $ >  >I:;9  (    :;9I  :;9   :;9I8  	I  
! I/  4 :;9I  .?:;9'I@�B  4 :;9I�B   I  .?:;9'@�B   :;9I   %�B   :;9I   I       '   I     	:;9  
 :;9I   :;9I  >I:;9  (   $ >  (    :;9I  :;9   :;9I8  $ >  I  ! I/  4 :;9I?<  !   >I:;9  ! I/  :;9   :;9I8  4 :;9I?<  :;9  4 G:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   :;9  & I  'I   I  '  I  ! I/  4 :;9I  4 :;9I  .?:;9'I@�B   :;9I  4 :;9I�B   :;9I�B  4 :;9I�B  4 :;9I  ��1  �� �B  ��1  1R�BXYW    1�B  !  "4 1�B  #1R�BUXYW  $U  %1R�BXYW  &�� 1  '.?:;9'I   ( :;9I  )4 :;9I  *.:;9'@�B  +.:;9'I   , :;9I  -.:;9'I@�B  ..:;9'   / :;9I  0.1@�B  14 1  21U  3�� �B1  4. ?<n:;9  5. ?<n:;   %�B   :;9I  $ >  $ >     >I:;9  (   (   	:;9  
 :;9I8   I  4 :;9I?<  :;9  I  ! I/   :;9I8   'I  '   I  'I  :;9   :;9I8       4 :;9I  4 G:;9  4 G:9  4 :;9I  4 :;9I?  4 :;9I  .?:;9'@�B    :;9I  !4 :;9I�B  "4 :;9I�B  #U  $1R�BUXYW  % 1�B  &U  '4 1�B  (1XYW  ) 1  *  +��1  ,�� �B  -��  .�� 1  /1R�BXYW  0.:;9'   1 :;9I  24 :;9I  3.:;9'I@�B  44 :;9I  5.:;9'I   6. ?:;9'@�B  7.?:;9'I@�B  8 :;9I�B  94 :;9I  :��1  ; :;9I  <1R�BUXYW  =���B1  >. :;9'   ?.?:;9'   @4 :;9I  A.:;9'I   B.:;9'I@�B  C4 :;9I�B  D.1@�B  E4 1  F  G4 1  H��  I.1@�B  J. ?<n:;9  K. ?<n:;   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  I  ! I/  (   :;9   :;9I8  :;9   :;9I8       ! I/  '   I  :;9   :;9I   :;9I  (    :;9I  :;9    :;9I8  !4 :;9I?<  "!   #>I:;9  $:;9  % '  &'I  ' :;9I8  (:;9  ):;9  * :;9I8  +4 G:;9  ,4 :;9I?  -4 G:;  .4 :;9I?  /4 :;9I  04 :;9I  1.?:;9'@�B  24 :;9I�B  3  44 :;9I�B  5�� 1  6��1  7�� �B  84 :;9I  9��1  :1R�BXYW  ; 1�B  <  =4 1  >1R�BUXYW  ?U  @4 1�B  A.:;9'   B���B1  C.?:;9'   D  E.:;9'I   F :;9I  GU  H 1R�BXYW  I. ?:;9'   J. ?:;9'I   K4 :;9I  L.?:;9'   M4 :;9I  N4 :;9I  O4 :;9I  P.?:;9'@�B  Q4 :;9I�B  R. 1@�B  S.1@�B  T�� �B1  U4 1  V. ?<n:;9  W. ?<n:;   %�B  $ >  $ >  >I:;9  (   (    :;9I  :;9  	 :;9I8  
 :;9I8  I  ! I/  4 :;9I  .?:;9'I@�B   :;9I�B   I   :;9I  4 :;9I�B  4 :;9I�B  ��1  �� �B   :;9I�B  .?:;9'I@�B   %�B   :;9I  $ >  $ >     :;9   :;9I8   I  	4 :;9I?<  
>I:;9  (   (   & I  (   :;9  I  ! I/   :;9I8       '   I  ! I/  :;9   :;9I   :;9I  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  " <  #:;9  $ :;9I8  %'I  &4 G:;9  '4 :;9I  (.?:;9'@�B  )1R�BUXYW  * 1�B  +��1  ,�� �B  -��1  .U  /4 1�B  0�� 1  1.:;9'   2 :;9I  34 :;9I  4.:;9'@�B  5 :;9I�B  64 :;9I�B  7 1  8�� �B1  94 :;9I  :. ?<n:;9  ;. ?<n:;   %�B  $ >   :;9I     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  :;9  I  ! I/  (   'I   I  '  ! I/       :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9   :;9I8   4 :;9I?<  !!   ">I:;9  #:;9  $ :;9I8  % :;9I8  &:;9  ' :;9I8  (4 :;9I?  )4 :;9I  *4 :;9I?  +.?:;9'@�B  ,1R�BUXYW  -U  .4 1�B  /�� �B1  0��1  1�� �B  2���B1  3.:;9'   44 :;9I  54 :;9I�B  64 :;9I�B  74 :;9I  8��1  9 :;9I  : :;9I�B  ; :;9I�B  <�� 1  =���B1  >.?:;9'I   ? :;9I  @.?:;9'   A4 :;9I  B
 :;9  C.?:;9'@�B  D4 :;9I�B  E4 :;9I�B  F4 :;9I  G.?:;9'I@�B  H :;9I�B  I  J4 :;9I  K.1@�B  L4 1  M4 1  N
 1  O 1�B  P1U  Q. ?<n:;9   %�B   :;9I  $ >  :;9   :;9I8   I  $ >  4 :;9I?<  	>I:;9  
(   (   I  ! I/  4 :;9I  4 :;9I  .?:;9'I@�B   :;9I�B   :;9I�B  4 :;9I�B  4 :;9I  ��  �� �B  ��1  ��  'I   I  .?:;9'I@�B   :;9I�B   :;9I�B  �� 1  ��1    :;9I  !4 :;9I�B  "4 :;9I�B  #.?:;9'@�B  $�� �B1  %. ?<n:;9   %U�B  $ >  $ >   :;9I     :;9   :;9I8   I  	4 :;9I?<  
>I:;9  (   (   & I  (   I  ! I/  :;9   :;9I8       ! I/  '   I  :;9   :;9I   :;9I  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  ":;9  # :;9I8  $ '  %'I  & :;9I8  ':;9  (:;9  ) :;9I8  *(   +4 :;9I?  ,4 G:;9  -4 G:;  .4 :;9I  /4 :;9I  04 :;9I?  1.?:;9'I@�B  24 :;9I�B  3  44 :;9I�B  5�� 1  6��1  7�� �B  8.?:;9'@�B  9 :;9I�B  :1R�BXYW  ; 1�B  <  =��1  >.:;9'I   ? :;9I  @4 :;9I  A :;9I  B :;9I�B  C4 1�B  D�� �B1  E���B1  F.:;9'   G4 :;9I  H :;9I  I.?:;9'   J. ?:;9'@�B  K4 :;9I  LU  M1  N  O1R�BUXYW  PU  Q4 1  R1R�BUXYW  S.:;9'I   T :;9I  U.?:;9'I@�B  V :;9I  W4 :;9I�B  X.1@�B  Y1U  Z. ?<n:;9  [. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  :;9  I  ! I/       '   I  :;9   :;9I   :;9I  ! I/   :;9I8  (    :;9I  :;9   :;9I8  4 :;9I?<  !    >I:;9  !:;9  " :;9I8  # :;9I8  $:;9  %:;9  & :;9I8  ':;9  ( :;9I8  ) '  *.?:;9'@�B  + :;9I�B  ,��1  -�� �B  .4 :;9I�B  /���B1  0.?:;9'I@�B  1��1  2 :;9I  31R�BUXYW  4 1�B  5 :;9I  61R�BUXYW  7.?:;9'@�B  8 :;9I�B  94 :;9I�B  : :;9I�B  ; :;9I  <1R�BXYW  = :;9I  > 1  ?4 :;9I�B  @�� 1  A�� �B1  B.?:;9'I@�B  C.?:;9'   D :;9I  E. ?:;9'@�B  F.1@�B  G 1  H. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  (   :;9  I  ! I/       '   I  :;9   :;9I   :;9I  ! I/   :;9I8  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  ":;9  # :;9I8  $:;9  % :;9I8  &'I  '4 G:;9  (4 :;9I?  )4 :;9I  *4 :;9I  +4 :;9I  ,.?:;9'I@�B  - :;9I�B  .4 :;9I�B  /4 :;9I�B  0��1  1�� �B  2�� 1  3��1  4.?:;9'@�B  5 :;9I  6���B1  74 :;9I  8 1R�BXYW  9. ?:;9'   :. 1@�B  ;. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
& I  I  ! I/  :;9  '   I  !   >I:;9  (        :;9   :;9I   :;9I  (    :;9I  :;9   :;9I8  ! I/  4 :;9I?<  >I:;9  (    4 G:;9  !4 G:;9   %�B   :;9I  $ >  :;9   :;9I8   I  $ >  4 :;9I?<  	4 G:;9  
.?:;9'I   :;9I  . ?:;9'I  .?:;9'I@�B   :;9I  .?:;9'I   . ?:;9'@�B  . ?:;9'I   . 1@�B  .1@�B   1   %�B   :;9I  $ >  :;9   :;9I8   I  $ >  4 :;9I?<  	>I:;9  
(   (   .?:;9'@�B   :;9I   %�B   :;9I  $ >  $ >  :;9   :;9I8   I  4 :;9I?<  	4 :;9I  
I  ! I/  .?:;9'@�B  4 :;9I�B  U  4 :;9I  ��1  �� �B  ��1  . ?:;9'  . ?:;9'   . ?:;9'  . 1@�B  . ?<n:;9   %�B   :;9I  $ >  :;9   :;9I8   I  $ >  4 :;9I?<  	>I:;9  
(   (   :;9  '   I  'I  4 :;9I  I  ! I/  4 :;9I?  4 :;9I?  .:;9'I    :;9I  4 :;9I  4 :;9I  .:;9'    :;9I  .:;9'@�B   :;9I�B   :;9I�B  4 :;9I   :;9I   4 :;9I�B  !.?:;9'@�B  "�� 1  #��1  $�� �B  %��1  &.:;9'I@�B  '4 :;9I�B  (1R�BUXYW  ) 1�B  *U  +4 1�B  ,.:;9'I@�B  - :;9I�B  . :;9I  /4 :;9I�B  04 :;9I�B  1.?:;9'@�B  2 :;9I  3.1@�B  44 1  51U  61UXYW  71R�BUXYW  8���B1  9. ?<n:;9  :. ?<n:;   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   I  ! I/  :;9  'I   I   '  '   'I  4 G:;9  4 :;9I  4 :;9I  . ?:;9'  . ?:;9'I@  . ?:;9'@  .?:;9'@�B   :;9I�B  ���B  �� �B  .?:;9'I@�B    :;9I�B  !. ?:;9'   ".:;9'   # :;9I  $. ?:;9'@  %.?:;9'@�B  & :;9I�B  '4 :;9I�B  (1R�BXYW  ) 1�B  *  +4 1�B  ,��1  -�� 1  ..:;9'   /4 :;9I  0 :;9I  1.:;9'I   2 :;9I  3. 1@�B  4. ?<n:;9   %�B   :;9I  $ >  $ >      I  I  ! I/  	:;  
 :;I8  :;9   :;9I8   I  4 :;9I?<  & I  >I:;9  (   (    '  :;9  'I   I  '  4 :;9I  4 :;9I  .?:;9'I@�B   :;9I�B    4 :;9I�B  4 :;9I  ��1   �� �B  !��1  ".?:;9'@�B  #   $4 :;9I�B  %1R�BXYW  & 1�B  '4 1  (4 1�B  )�� 1  *! I/  +.:;9'I   , :;9I  -4 :;9I  .4 :;9I  /. :;9'I   0.?:;9'@�B  14 :;9I�B  2. ?:;9'I   3.?:;9'@�B  4 :;9I�B  5�� �B1  64 :;9I�B  7���B1  8 :;9I�B  9.?:;9'I@�B  :4 :;9I  ;1R�BXYW  < 1  =.:;9'I   > :;9I  ? :;9I  @ :;9I  A. 1@�B  B. ?<n:;9  C. ?<n:;   %�B  $ >   :;9I  $ >  4 :;9I?<   I  4 :;9I  . ?:;9'@�B  	.?:;9'@�B  
 :;9I   :;9I�B  ���B1  �� �B  .?:;9'I@�B  4 :;9I�B  1R�BUXYW  �� 1  . ?:;9'I   .1@�B  �� �B1  . ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
 :;9I8  >I:;9  (   .?:;9'I@�B   :;9I�B  4 :;9I�B  ��1  �� �B   :;9I  .?:;9'@�B  �� 1  ���B1   :;9I   :;9I�B    ��1  &   . ?<n:;9  . ?<n:;   %�B   :;9I  $ >  :;9   :;9I8   I  $ >  4 :;9I?<  	>I:;9  
(   (   4 G:;9  .?:;9'I@�B  4 :;9I�B  ��1  �� �B  .?:;9'@�B  4 :;9I  .:;9'    :;9I   :;9I�B  ���B1  . ?<n:;9   %�B   :;9I  $ >  >I:;9  (   $ >  .?:;9'@�B   :;9I  	 I  
.?:;9'@�B   %�B   :;9I  $ >  $ >  >I:;9  (   (   :;9  	 :;9I8  
I  ! I/  .?:;9'@�B   :;9I�B   :;9I�B   I  .?:;9'I@�B   :;9I   %�B   :;9I  $ >     :;9   :;9I8   I  & I  	$ >  
4 :;9I?<  >I:;9  (   (   4 :;9I?  4 :;9I  :;9  I  ! I/  4 :;9I  .?:;9'I@�B   :;9I�B  4 :;9I�B  ���B1  �� �B  ��1  ��1  .?:;9'@�B   :;9I�B  1R�BXYW    4 1�B   �� �B1  !.:;9'I   "4 :;9I  #1R�BUXYW  $ 1�B  %U  &.:;9'I@�B  '4 :;9I�B  ( :;9I  ). ?:;9'   *.:;9'   + :;9I  , :;9I  -.1@�B  .4 1  /1  0�� 1  1. 1@�B  2. ?<n:;9   %�B   :;9I  $ >  :;9   :;9I8   I  $ >  4 :;9I?<  	4 :;9I?  
I  ! I/  . ?:;9'@�B  .?:;9'@�B   :;9I�B  4 :;9I  4 :;9I�B  ��1  �� �B  ��1  ���B1  .?:;9'@�B  . ?<n:;9   %�B  $ >  $ >   :;9I  .?:;9'I@�B   :;9I   :;9I�B    	4 :;9I�B  
.?:;9'I@�B   %U�B   :;9I  $ >  $ >     :;9   :;9I8   I  	4 :;9I?<  
>I:;9  (   (   & I  (   I  !   :;9   '  ! I/  'I   I  '  ! I/       :;9   :;9I   :;9I   :;9I8  (    :;9I   :;9  ! :;9I8  "4 :;9I?<  #>I:;9  $:;9  % :;9I8  & :;9I8  ':;9  (:;9  ) :;9I8  *4 G:;9  +4 :;9I?  ,(   -4 :;9I?  .4 :;9I?  /4 :;9I  0. ?:;9'@�B  1.?:;9'@�B  2 :;9I  3. ?:;9'   4.?:;9'@�B  54 :;9I  64 :;9I�B  74 :;9I�B  8U  9��1  :�� �B  ;��1  <�� 1  =.?:;9'I@�B  > :;9I�B  ? 1R�BXYW  @1R�BXYW  A 1�B  B��  C.:;9'I   D :;9I  E :;9I�B  F.?:;9'I@�B  G�� �B1  H���B1  I.?:;9'   J :;9I  K1R�BUXYW  LU  M4 1�B  N4 :;9I  O1R�BXYW  P 1R�BUXYW  Q4 :;9I  R.1@�B  S1  T1U  U1  V4 1  W. 1@�B  X���B1  Y. ?<n:;9  Z. ?<n:;   %�B   :;9I  $ >   I  I  ! I/  :;   :;I8  	   
:;9   :;9I8   I  & I  $ >  4 :;9I?<  >I:;9  (   (   :;9  'I   I  '  .?:;9'I@�B   :;9I�B   :;9I�B     4 :;9I  4 :;9I�B  ��1  �� �B  .?:;9'I     :;9I  ! :;9I  "4 :;9I  #4 :;9I  $��1  %���B1  &4 :;9I�B  '.?:;9'@�B  ( :;9I�B  )4 :;9I�B  *�� 1  +4 :;9I�B  ,.?:;9'I@�B  - :;9I�B  .4 :;9I  /.1@�B  0 1�B  14 1  21U  3 1  4U  54 1�B  6. ?<n:;9   %�B  I  ! I/  & I  $ >  4 :;9I  4 :;9I?  $ >  	. ?:;9'@�B  
. ?:;9'I@�B   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  (   I  ! I/  ! I/       '   I  :;9   :;9I   :;9I  :;9   :;9I8  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  ":;9  # :;9I8  $ :;9I8  %:;9  &:;9  ' :;9I8  ( '  )(   *4 G:;9  +.?:;9'I@�B  , :;9I  -4 :;9I�B  ..?:;9'@�B  / :;9I�B  0��1  1�� �B  2.?:;9'@�B  3 :;9I  44 :;9I�B  5.?:;9'I@�B  6 :;9I�B  74 :;9I�B  8��1  9���B1  :. ?<n:;9  ;. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  (   I  ! I/  ! I/       '   I  :;9   :;9I   :;9I  :;9   :;9I8  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  ":;9  # :;9I8  $ :;9I8  %:;9  &:;9  ' :;9I8  ( '  )(   *.?:;9'@�B  + :;9I�B  , :;9I�B  -4 :;9I�B  .��1  /�� �B  0��1  14 :;9I�B  24 :;9I  3  4���B1  5�� 1  6.?:;9'I@�B  7 :;9I�B  84 :;9I�B  9�� �B1  :.?:;9'@�B  ;���B1  <. ?<n:;9  =. ?<n:;  >. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  :;9   '  (   I  ! I/  ! I/       '   I  :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9   :;9I8   4 :;9I?<  !!   ">I:;9  #:;9  $ :;9I8  % :;9I8  &:;9  ':;9  ( :;9I8  )(   *4 :;9I?  +4 :;9I?  ,.?:;9'@�B  - :;9I�B  .4 :;9I�B  /�� �B1  0.?:;9'   1 :;9I  24 :;9I  34 :;9I  4��1  5�� �B  6���B1  74 :;9I  84 :;9I�B  9�� 1  : :;9I�B  ;1R�BUXYW  < 1�B  =.:;9'I   > :;9I  ?.?:;9'I   @��1  A���B1  B
 :;9  C  D1R�BXYW  E.?:;9'I@�B  F.?:;9'I   G :;9I  H4 :;9I  I4 :;9I  J.?:;9'@�B  K :;9I�B  L.?:;9'   M :;9I  N.1@�B  O4 1  P1U  QU  R4 1�B  S1  T  U1  V 1  W. ?<n:;9  X. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  (   I  ! I/  ! I/       '   I  :;9   :;9I   :;9I  :;9   :;9I8  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  ":;9  # :;9I8  $ :;9I8  %:;9  &:;9  ' :;9I8  ( '  )(   *.?:;9'I@�B  + :;9I�B  ,4 :;9I�B  -4 :;9I�B  .��1  /�� �B  0��1  1.?:;9'I@�B  2 :;9I�B  34 :;9I�B  4  5.?:;9'   6 :;9I  74 :;9I  8.1@�B  9 1�B  :4 1�B  ;1U  <U  =4 1  >���B1  ?. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  (   (   I  !   ! I/  :;9   '  '   I   :;9I8       ! I/  :;9   :;9I   :;9I   :;9I  :;9    :;9I8  !4 :;9I?<  ">I:;9  #:;9  $ :;9I8  % :;9I8  &:;9  ':;9  ( :;9I8  )(   *4 G:;9  +.?:;9'@�B  , :;9I�B  -4 :;9I�B  .4 :;9I�B  /�� 1  0��1  1�� �B  2���B1  3���B1  4��1  51R�BUXYW  6 1�B  7 1  8U  94 1�B  :1R�BXYW  ;1U  <.?:;9'I   = :;9I  > :;9I  ?.?:;9'I   @ :;9I  A4 :;9I  B.?:;9'I@�B  C :;9I  D :;9I�B  E :;9I�B  F4 :;9I�B  G :;9I  H.1@�B  I1U  J4 1  K 1  L1  M. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  I  ! I/  ! I/       '   I  :;9   :;9I   :;9I  :;9   :;9I8  (    :;9I  :;9   :;9I8  4 :;9I?<  !    >I:;9  !:;9  " :;9I8  # :;9I8  $:;9  %:;9  & :;9I8  ' '  ((   ).?:;9'@�B  * :;9I�B  +4 :;9I�B  ,��1  -�� �B  .��1  /.?:;9'   0 :;9I  14 :;9I�B  2.?:;9'@�B  3 :;9I�B  44 :;9I�B  54 :;9I�B  6�� 1  7.?:;9'   8 :;9I  94 :;9I  :.1@�B  ; 1  <1  = 1�B  >4 1  ?  @4 1�B  A1U  B. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
& I  >I:;9  (   (   :;9   '  (   I  ! I/  ! I/       '   I  :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9   :;9I8   4 :;9I?<  !!   ">I:;9  #:;9  $ :;9I8  % :;9I8  &:;9  ':;9  ( :;9I8  )(   *4 :;9I?  +4 :;9I?  ,4 G:;9  -4 :;9I?  .4 G:;9  /.:;9'   0 :;9I  14 :;9I  24 :;9I  3  44 :;9I  5.?:;9'I@�B  6 :;9I�B  74 :;9I�B  8��1  9�� �B  :.?:;9'I   ; :;9I  <.?:;9'@�B  =4 :;9I�B  >���B1  ? :;9I�B  @��1  A
 :;9  B�� 1  C���B1  D.?:;9'   E.?:;9'I   F :;9I  G.?:;9'I@�B  H :;9I�B  I :;9I�B  J4 :;9I�B  K4 :;9I�B  L :;9I  M4 :;9I  N.1@�B  O 1�B  P4 1  Q1U  RU  S4 1�B  T1  U1R�BXYW  V  W. ?<n:;9  X. ?<n:;9   %�B   :;9I  $ >  $ >     & I  >I:;9  (   	:;9  
 :;9I8   I  4 :;9I?<  (   (   I  ! I/  :;9   :;9I8       ! I/  '   I  :;9   :;9I   :;9I  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  ":;9  # :;9I8  $ :;9I8  %:;9  &:;9  ' :;9I8  ( '  )'I  *(   +4 G:;9  ,4 :;9I?  -4 :;9I  ..?:;9'I@�B  / :;9I�B  0 :;9I�B  14 :;9I�B  24 :;9I�B  3��1  4�� �B  5�� 1  6���B1  7.:;9'   8 :;9I  94 :;9I  :.:;9'@�B  ;��  <4 :;9I  =1R�BXYW  > 1�B  ?  @4 1  A��1  B.?:;9'I@�B  C.?:;9'@�B  D :;9I  E.?:;9'I@�B  F :;9I�B  G4 :;9I  H4 :;9I�B  I�� �B1  J.?:;9'@�B  K :;9I  L :;9I�B  M4 :;9I�B  N.?:;9'I   O :;9I  P :;9I  Q4 :;9I  R4 :;9I  S.1@�B  T4 1�B  U1  V. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  :;9   '  (   I  ! I/  ! I/       '   I  :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9   :;9I8   4 :;9I?<  !!   ">I:;9  #:;9  $ :;9I8  % :;9I8  &:;9  ':;9  ( :;9I8  )(   *4 :;9I?  +4 G:;9  ,.?:;9'@�B  - :;9I�B  .4 :;9I�B  /4 :;9I�B  0��1  1�� �B  2�� 1  3�� �B1  4.?:;9'I@�B  5��1  6  74 :;9I  8 :;9I�B  9���B1  :���B1  ;4 :;9I  <4 :;9I  =.?:;9'@�B  > :;9I�B  ?4 :;9I�B  @U  A.?:;9'   B :;9I  C4 :;9I  D.?:;9'I@�B  E :;9I�B  F4 :;9I�B  G��  H.1@�B  I 1�B  J4 1  K1U  LU  M4 1�B  N. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  :;9   '  (   I  ! I/  ! I/       '   I  :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9   :;9I8   4 :;9I?<  !!   ">I:;9  #:;9  $ :;9I8  % :;9I8  &:;9  ':;9  ( :;9I8  )(   *4 G:;9  +.?:;9'@�B  , :;9I�B  -4 :;9I�B  .��1  /�� �B  0���B1  1 :;9I  2.?:;9'@�B  3 :;9I  44 :;9I�B  5.?:;9'I@�B  6 :;9I�B  74 :;9I�B  8�� 1  9���B1  :�� �B1  ;. ?<n:;9  <. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  (   I  ! I/  ! I/       '   I  :;9   :;9I   :;9I  :;9   :;9I8  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  ":;9  # :;9I8  $ :;9I8  %:;9  &:;9  ' :;9I8  ( '  )(   *4 :;9I?  +4 :;9I?  ,.?:;9'@�B  - :;9I�B  .4 :;9I�B  /4 :;9I�B  0��1  1�� �B  2���B1  3 :;9I�B  4��1  5�� 1  6 :;9I  7 :;9I  8�� �B1  9.:;9'@�B  :���B1  ;4 :;9I  <.?:;9'   = :;9I  >4 :;9I  ?.?:;9'I   @.?:;9'@�B  A :;9I�B  B4 :;9I�B  C4 :;9I�B  D��  E.1@�B  F 1�B  G4 1�B  H1U  I 1  JU  K4 1  L1U  M. ?<n:;9  N. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
I  !   >I:;9  (   (   & I  :;9   '  ! I/  ! I/  (        '   I  :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9    :;9I8  !4 :;9I?<  ">I:;9  #:;9  $ :;9I8  % :;9I8  &:;9  ':;9  ( :;9I8  )(   *4 G:;9  +4 :;9I?  ,4 :;9I?  -.?:;9'@�B  .4 :;9I�B  /1R�BUXYW  0 1�B  1U  24 1�B  3��1  4�� �B  5�� 1  6��1  74 :;9I�B  81R�BXYW  9���B1  :���B1  ;4 :;9I  < 1  =  >.?:;9'I@�B  ?4 :;9I  @ :;9I�B  A.:;9'   B :;9I  C4 :;9I  D.:;9'@�B  E :;9I�B  F�� �B1  G1R�BUXYW  H1R�BXYW  I1R�BXYW  J.:;9'   K :;9I  L. :;9'I   M.:;9'@�B  N4 :;9I�B  O4 :;9I�B  P :;9I�B  Q.:;9'I@�B  R :;9I  S.:;9'I   T4 :;9I  U.?:;9'I@�B  V4 :;9I  W.1@�B  X1  Y4 1  Z  [4 1  \. ?<n:;9  ]. ?<n:;9  ^. ?<n:;   %�B  $ >   :;9I     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  (   :;9   '  'I   I  '  I  ! I/  ! I/       :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9    :;9I8  !4 :;9I?<  "!   #>I:;9  $:;9  % :;9I8  & :;9I8  ':;9  (:;9  ) :;9I8  *(   +4 G:;9  ,4 :;9I  -.?:;9'@�B  .�� 1  /�� �B1  0 :;9I�B  1 :;9I�B  24 :;9I�B  34 :;9I  44 :;9I�B  51R�BXYW  6 1�B  7  84 1�B  91R�BUXYW  :U  ;4 1  <��1  =�� �B  >��1  ?.:;9'   @ :;9I  A4 :;9I  B :;9I  C4 :;9I  D4 :;9I  E���B1  F.?:;9'@�B  G :;9I�B  H4 :;9I�B  I4 :;9I�B  J4 :;9I  K.?:;9'I   L.1@�B  M. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  :;9   '  I  ! I/  ! I/       '   I  :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  ":;9  # :;9I8  $ :;9I8  %:;9  &:;9  ' :;9I8  ((   )4 :;9I?  *4 :;9I?  +.?:;9'I@�B  , :;9I�B  -4 :;9I�B  .4 :;9I�B  /�� �B1  0 :;9I�B  1��1  2�� �B  3�� 1  4��1  5.?:;9'I@�B  6 :;9I�B  74 :;9I�B  84 :;9I�B  94 :;9I  :.?:;9'I   ; :;9I  < :;9I  =4 :;9I  >4 :;9I  ?.1@�B  @ 1�B  A 1  B4 1�B  C1U  DU  E4 1  F. ?<n:;9   %�B   :;9I  $ >  $ >     :;9   :;9I8   I  	4 :;9I?<  
>I:;9  (   (   & I  (   I  ! I/  :;9   :;9I8       ! I/  '   I  :;9   :;9I   :;9I  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  ":;9  # :;9I8  $ '  %'I  & :;9I8  ':;9  (:;9  ) :;9I8  *(   +4 :;9I?  ,4 G;9  -4 G:;9  .4 G;9  /.?:;9'@�B  04 :;9I�B  14 :;9I�B  2��1  3�� �B  4��1  5.?:;9'I@�B  6 :;9I�B  71R�BXYW  8 1�B  9  :4 1<  ;1  <4 1�B  =.:;9'   > :;9I  ?4 :;9I  @  A4 :;9I  B�� 1  C�� �B1  D���B1  E :;9I�B  F :;9I  G.?:;9'I@�B  H :;9I  I :;9I  J :;9I�B  K.?:;9'@�B  L4 :;9I  M4 :;9I�B  N. ?<n:;9  O. ?<n:;9  P. ?<n:;   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  :;9   '  (   I  ! I/  ! I/       '   I  :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9   :;9I8   4 :;9I?<  !!   ">I:;9  #:;9  $ :;9I8  % :;9I8  &:;9  ':;9  ( :;9I8  )(   *4 :;9I?  +4 G:;  ,.?:;9'I@�B  - :;9I�B  .��1  /�� �B  0�� 1  1��1  2.?:;9'@�B  3 :;9I�B  44 :;9I�B  54 :;9I�B  6���B1  7.?:;9'   8 :;9I  9 :;9I  :4 :;9I  ;.1@�B  < 1�B  =4 1�B  >1  ? 1  @  A. ?<n:;9  B. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  (   I  ! I/  :;9   :;9I8       ! I/  '   I  :;9   :;9I   :;9I  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  ":;9  # :;9I8  $ '  % :;9I8  &:;9  ':;9  ( :;9I8  )(   *.?:;9'I@�B  + :;9I�B  ,4 :;9I�B  -4 :;9I�B  .��1  /�� �B  0��1  1. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  I  ! I/  ! I/  (        '   I  :;9   :;9I   :;9I  :;9   :;9I8  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  ":;9  # :;9I8  $ :;9I8  %:;9  &:;9  ' :;9I8  ( '  )(   *4 G:;9  +.?:;9'@�B  ,4 :;9I�B  -�� 1  .4 :;9I�B  /��1  0�� �B  1��  2 :;9I  3. ?:;9'@�B  4. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  (   I  ! I/  ! I/       '   I  :;9   :;9I   :;9I  :;9   :;9I8  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  ":;9  # :;9I8  $ :;9I8  %:;9  &:;9  ' :;9I8  ( '  )(   *4 :;9I?  +.?:;9'@�B  , :;9I�B  -4 :;9I�B  .4 :;9I�B  /���B1  0�� �B  1�� 1  2��1  3��1  4���B1  5.?:;9'   6 :;9I  74 :;9I  84 :;9I  9.1@�B  : 1�B  ;4 1  <1  =  >4 1�B  ?. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  (   :;9   '  I  ! I/  ! I/       '   I  :;9   :;9I   :;9I  (    :;9I  :;9   :;9I8  4 :;9I?<   !   !>I:;9  " :;9I8  #:;9  $ :;9I8  % :;9I8  &:;9  ':;9  ( :;9I8  )4 :;9I?  *4 :;9I?  +.?:;9'@�B  , :;9I�B  -4 :;9I�B  .4 :;9I�B  /�� �B1  0��1  1�� �B  2�� 1  3��1  4 :;9I�B  5.?:;9'I@�B  64 :;9I  7.?:;9'@�B  8 :;9I�B  94 :;9I�B  :
 :;9  ;. ?:;9'@�B  <4 :;9I�B  =���B1  >
 :;9  ?. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  :;9   '  (   'I   I  '  I  ! I/  ! I/       :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9    :;9I8  !4 :;9I?<  "!   #>I:;9  $:;9  % :;9I8  & :;9I8  ':;9  (:;9  ) :;9I8  *(   +4 G:;9  ,4 :;9I?  -4 :;9I?  ..?:;9'@�B  /4 :;9I�B  04 :;9I�B  14 :;9I  2��1  3�� �B  4�� �B1  5.?:;9'I@�B  6 :;9I�B  7��1  8.?:;9'I   9 :;9I  :4 :;9I  ;4 :;9I  <�� 1  =1R�BXYW  >  ?4 1�B  @.:;9'   A :;9I�B  B.?:;9'@�B  C :;9I�B  D4 :;9I�B  E4 :;9I�B  F4 :;9I  G���B1  H :;9I  I.1@�B  J 1�B  K4 1  L1U  MU  N. ?<n:;9  O. ?<n:;   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  (   :;9   '  'I   I  '  I  ! I/  ! I/       :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9    :;9I8  !4 :;9I?<  "!   #>I:;9  $:;9  % :;9I8  & :;9I8  ':;9  (:;9  ) :;9I8  *4 :;9I?  +4 G:;9  ,4 :;9I  -4 :;9I?  .4 G:;9  /.?:;9'@�B  04 :;9I�B  14 :;9I�B  2��1  3�� �B  4���B1  5 :;9I�B  6 :;9I�B  74 :;9I  8�� 1  9�� �B1  : :;9I  ;��1  <4 :;9I  =.?:;9'@�B  >4 :;9I�B  ?4 :;9I�B  @. ?<n:;9   %�B   :;9I  $ >  $ >     :;9   :;9I8   I  	4 :;9I?<  
>I:;9  (   (   & I  :;9       I  ! I/  ! I/  '   I  :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9   :;9I8  4 :;9I?<  !    >I:;9  !:;9  " :;9I8  # :;9I8  $:;9  %:;9  & :;9I8  ' '  (4 :;9I?  )4 G:;9  *4 :;9I?  +.?:;9'@�B  , :;9I�B  -��1  .�� �B  /�� 1  0�� �B1  1 :;9I  24 :;9I�B  3.?:;9'I@�B  4 :;9I�B  54 :;9I�B  6��1  71R�BXYW  8 1  94 :;9I  :.?:;9'   ; :;9I  <. ?:;9'   =���B1  >.?:;9'I@�B  ? :;9I�B  @ :;9I�B  A4 :;9I�B  B4 :;9I�B  C.?:;9'@�B  D :;9I  E. 1@�B  F.1@�B  G 1  H. ?<n:;9  I. ?<n:;   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  :;9   '  (   'I   I  '  I  ! I/   :;9I8       ! I/  :;9   :;9I   :;9I  (    :;9I  :;9    :;9I8  !4 :;9I?<  "!   #>I:;9  $:;9  % :;9I8  & :;9I8  ':;9  (:;9  ) :;9I8  *4 G:;9  +4 :;9I?  ,.?:;9'@�B  -4 :;9I�B  .4 :;9I�B  /��1  0�� �B  1�� 1  2��1  3.?:;9'@�B  4 :;9I�B  5.?:;9'I@�B  6 :;9I  7 :;9I�B  8.?:;9'I@�B  9 :;9I�B  :4 :;9I�B  ;.?:;9'@�B  <4 :;9I�B  =.?:;9'@  > :;9I�B  ?. ?:;9'@�B  @. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  :;9   '  (   I  ! I/   :;9I8       ! I/  '   I  :;9   :;9I   :;9I  (    :;9I  :;9   :;9I8   4 :;9I?<  !!   ">I:;9  #:;9  $ :;9I8  % :;9I8  &:;9  ':;9  ( :;9I8  )4 G:;9  *4 :;9I?  +.?:;9'@�B  , :;9I�B  -4 :;9I�B  .4 :;9I  /4 :;9I�B  0��1  1�� �B  2�� 1  3.?:;9'@�B  44 :;9I  54 :;9I�B  64 :;9I�B  7��1  8.?:;9'@�B  9 :;9I�B  :. ?<n:;9   %�B   :;9I  & I  $ >  $ >     :;9   :;9I8  	 I  
4 :;9I?<  >I:;9  (   (        '   I  :;9   :;9I   :;9I  I  ! I/  ! I/  :;9   :;9I8  (    :;9I  :;9   :;9I8  4 :;9I?<  !    >I:;9  !:;9  " :;9I8  # :;9I8  $:;9  % :;9I8  &4 :;9I?  '4 G:;9  (. ?:;9'@�B   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  (   :;9   '  'I   I  '  I  ! I/  ! I/       :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9    :;9I8  !4 :;9I?<  "!   #>I:;9  $:;9  % :;9I8  & :;9I8  ':;9  (:;9  ) :;9I8  *4 G:;9  +4 :;9I?  ,4 G:;9  -4 :;9I?  .4 :;9I  /.?:;9'@�B  04 :;9I�B  1�� 1  2��1  3�� �B  4�� �B1  5 :;9I�B  64 :;9I�B  7���B1  8��1  9 :;9I�B  :.?:;9'@�B  ;. ?:;9'I@�B  <. ?:;9'@�B  =.?:;9'@�B  > :;9I�B  ?4 :;9I�B  @4 :;9I�B  A. ?<n:;9   %�B   :;9I  $ >  :;9   :;9I8   I  $ >  4 :;9I?<  	 :;9I8  
I  ! I/  .?:;9'@�B   :;9I�B   :;9I�B  ���B1  �� �B  4 :;9I  ��1  .?:;9'@�B   :;9I�B   :;9I�B  4 :;9I�B  ��1  .:;9'@�B  4 :;9I    .?:;9'@�B   :;9I   %�B  $ >  $ >      :;9I  :;9   :;9I8   I  	I  
! I/  :;9  4 :;9I?<  !   >I:;9  (   4 G:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	& I  
4 :;9I?<  >I:;9  (   (   :;9  I  ! I/  ! I/       '   I  :;9   :;9I   :;9I  (    :;9I  :;9   :;9I8  4 :;9I?<  !    :;9I8   4 :;9I
  !4 :;9I  ". ?:;9'@�B  #.?:;9'@�B  $ :;9I�B  %��1  &�� �B  '. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  :;9  I  ! I/   '  'I   I  '       :;9   :;9I   :;9I  ! I/   :;9I8  (    :;9I  :;9   :;9I8   4 :;9I?<  !!   ">I:;9  #:;9  $ :;9I8  % :;9I8  &:;9  ':;9  ( :;9I8  )4 :;9I?  *.?:;9'@�B  + :;9I�B  , :;9I�B  -4 :;9I�B  .��1  /�� �B  0�� 1  1��1  2 :;9I  3 :;9I�B  4 :;9I�B  54 :;9I�B  6 :;9I  7���B1  81R�BUXYW  9 1�B  :4 :;9I  ;�� �B1  <.?:;9'   = :;9I  > :;9I  ?.1@�B  @ 1  A. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  :;9   '  (   'I   I  '  I  ! I/       :;9   :;9I   :;9I  ! I/   :;9I8  (    :;9I  :;9    :;9I8  !4 :;9I?<  "!   #>I:;9  $:;9  % :;9I8  & :;9I8  ':;9  (:;9  ) :;9I8  *(   +4 G:;9  ,4 :;9I  -4 :;9I  ..?:;9'@�B  /�� 1  0��1  1�� �B  2. ?:;9'   34 :;9I�B  4��1  5�� �B1  6���B1  7.:;9'@�B  8 :;9I�B  94 :;9I�B  :��  ;��  <4 :;9I  =.?:;9'I@�B  > :;9I�B  ?  @4 :;9I  A.1@�B  B. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  I  ! I/  :;9   '  '   I  (    :;9I8       ! I/  :;9   :;9I   :;9I  (    :;9I  :;9   :;9I8   4 :;9I?<  !!   ">I:;9  #:;9  $ :;9I8  % :;9I8  &:;9  ':;9  ( :;9I8  )(   *'I  +4 :;9I  ,4 G:;9  -.?:;9'@�B  .�� 1  /.?:;9'I@�B  0�� �B1  1 :;9I�B  24 :;9I�B  34 :;9I  4��1  5�� �B  6��1  7���B1  84 :;9I  94 :;9I�B  :4 :;9I  ;1R�BUXYW  < 1  = 1�B  >U  ?4 1�B  @.:;9'I@�B  A :;9I�B  B.:;9'I   C :;9I  D4 :;9I  E.?:;9'@�B  F :;9I�B  G4 :;9I�B  H  I.:;9'@�B  J4 :;9I�B  K. ?<n:;9   %�B  $ >   :;9I  $ >  & I  I  ! I/  4 :;9I?<  	 I  
! I/  4 G:;9  4 G:;9  .?:;9'I@�B   :;9I�B  4 :;9I�B   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   :;9  I  ! I/  'I   I  '  4 G:;9  4 :;9I?  4 :;9I  :;9   :;9I8   :;9I  .?:;9'@�B   :;9I�B  4 :;9I?<  4 :;9I�B  4 :;9I�B  ��1  �� �B   �� 1  !���B1  "4 :;9I  #4 :;9I  $��1  %�� �B1  &. ?:;9'@�B  ' :;9I  ( :;9I�B  ) :;9I  *��  +.?:;9'@�B  , :;9I�B  - :;9I�B  .4 :;9I�B  /4 :;9I�B  0��  1 :;9I  2.?:;9'   3 :;9I  4 :;9I  5.1@�B  6 1�B  71U  8 1  9. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (   (   & I  :;9   '  (   'I   I  '  I  ! I/  ! I/       :;9   :;9I   :;9I   :;9I8  (    :;9I  :;9    :;9I8  !4 :;9I?<  "!   #>I:;9  $:;9  % :;9I8  & :;9I8  ':;9  (:;9  ) :;9I8  *4 :;9I  +4 :;9I  ,4 :;9I  -4 :;9I  ..?:;9'@�B  / :;9I�B  0��1  1�� �B  2�� 1  3�� �B1  4.?:;9'   5 :;9I  6���B1  7.:;9'@�B  8��1  9.:;9'@�B  :4 :;9I�B  ;��  <��  =4 :;9I�B  >4 :;9I  ?.?:;9'I@�B  @ :;9I  A. ?:;9'@�B  B. ?:;9'<  C :;9I  D :;9I�B  E4 :;9I  F���B1  G  H :;9I  I.1@�B  J4 1  K  L4 1�B  M 1�B  N1U  O1U  P 1  QU  R 1  S1  T. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
 :;9I8  I  ! I/  :;9  'I   I  '  4 :;9I  .?:;9'@�B   :;9I�B  4 :;9I�B  1R�BUXYW   1�B  U  4 1  1R�BXYW    4 1�B  4 1  ��1  �� �B  ��1   .:;9'   ! :;9I  "4 :;9I  #.:;9'I   $4 :;9I  %. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
:;9  'I   I  '  I  ! I/  4 :;9I  .?:;9'I@�B   :;9I�B   :;9I�B  ���B  �� �B  .?:;9'@�B  4 :;9I  4 :;9I  ��1  . ?<n:;9   %�B   :;9I  $ >  $ >  >I:;9  (   (    I  	4 :;9I?<  
   :;9   :;9I8  :;9  'I   I  '  I  ! I/  .?:;9'I@�B  4 :;9I�B  4 :;9I�B    �� 1  ��1  �� �B  ��1  . ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  & I  	$ >  
4 :;9I?<  >I:;9  (   (   :;9  'I   I  '  I  ! I/  4 G:;9  4 :;9I  :;9   :;9I8  4 :;9I  .?:;9'@�B   :;9I�B  4 :;9I�B  4 :;9I�B  ��1  �� �B  ��1     !�� 1  "�� �B1  #���B1  $.?:;9'I@�B  % :;9I�B  &.?:;9I<  '   (.?:;9'I   ) :;9I  *4 :;9I  +4 :;9I  ,  -. ?:;9'I@�B  ..?:;9'I@�B  / :;9I�B  04 :;9I�B  14 :;9I�B  21R�BUXYW  3 1�B  4U  54 1�B  61  7.:;9'   8 :;9I  94 :;9I  :4 :;9I  ; :;9I�B  <.1@�B  =4 1  >1  ?  @. ?<n:;9  A. ?<n:;9   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
>I:;9  (    :;9I8  :;9  4 :;9I?  . ?:;9'I@�B  .?:;9'I@�B  4 :;9I�B  .?:;9'@�B   :;9I�B   :;9I�B  ��1  �� �B  ��1  �� 1  .?:;9'I@�B   :;9I�B   :;9I�B  4 :;9I�B  .?:;9'@�B  4 :;9I   :;9I   . ?<n:;9  !. ?<n:;   %�B   :;9I  $ >     :;9   :;9I8   I  $ >  	4 :;9I?<  
:;9  'I   I  '  >I:;9  (    :;9I8  4 G;9  .?:;9'I@�B   :;9I�B   :;9I�B  4 :;9I�B  4 :;9I  ��1  �� �B  ���B1  .:;9'@�B  �� 1  .:;9'I@�B  ��1  . ?<n:;9   %�B   :;9I  $ >  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<  >I:;9  (   (   :;9  '   I  'I  I  ! I/  ! I/  4 G:;9  4 :;9I  4 :;9I
  . ?:;9'@�B  .?:;9'@�B  4 :;9I  4 :;9I  1R�BUXYW   1�B  U  4 1�B   ��1  !�� �B  "��1  #.:;9'   $ :;9I  % :;9I  &4 :;9I  '.:;9'I   ( :;9I  ). ?<n:;9   %�B  I  ! I/  & I  $ >  4 :;9I   :;9I  $ >  	>I:;9  
(   (   4 :;9I?<   I  :;9   :;9I8   'I  ! I/   :;9I8  4 :;9I  4 :;9I?   :;9I8  4 G:;9  :;9  4 :;9I  . ?:;9'  .?:;9'@�B   :;9I  . ?:;9'    :;9I�B  ���B1  �� �B   .?:;9'I@�B  ! :;9I�B  "4 :;9I�B  #4 :;9I  $4 :;9I�B  %��1  &  '�� �B1  (. ?:;9'  ).?:;9'@�B  *�� 1  +4 :;9I�B  ,. ?:;9'I<  -��1  . :;9I�B  / :;9I  0. 1@�B  1. ?<n:;9  2. ?<n:;   %�B  $ >   :;9I  $ >  4 :;9I?<   I  4 G:;9  .?:;9@�B  	.?:;'I<  
 I  ��1  �� �B  �� �B1     . ?<n:;  . ?<n:;9   %U�B   :;9I  $ >     :;9   :;9I8   I  & I  	$ >  
4 :;9I?<   :;9I8  ;   9:;  9 :;9�  : :;9   :;9  .?:;9nI<   I  .?:;9nI<  9:;9  :;9n  .?:;9I<     &   I  .?:;9I<  .?:;9<  .?:;9�<  . ?:;9I<  :;9  .?:;9n2<d    I4  !.?:;9nI2<d  " :;9I82  # :;9I82  $/ I  % <  &  '.?n4<d  (I  )! I/  *4 :;9I  +4 :;9I?  ,.4@�B  -1R�BXYW  . 1�B  / 1  0.4   1 :;9I  2.?:;9@�B  3 :;9I�B  4��1  5�� �B  6�� �B1  7.?:;9I@�B  8 :;9I  9  :4 :;9I�B  ;4 :;9I  < :;9I�B  =�� 1  >��1  ?.:;9@�B  @4 :;9I�B  A1R�BUXYW  B.:;9I   C :;9I  D.G:;9d   E I4  F.1nd  G 1  H. ?<n:;9   %  $ >   :;9I  $ >  :;9n   :;9I8   :;9I8  .?:;9n@�B  	 :;9I  
4 :;9I  4 :;9I  .?:;9nI@�B   I   %   :;9I  $ >  $ >  :;9   :;9I8   :;9I8   I  	:;9n  
I  ! I/  & I  9:;  9 :;9�  : :;9   :;9  .?:;9nI<   I  .?:;9nI<  9:;9     .?:;9I<     &   I  .?:;9I<  .?:;9<  .?:;9�<  . ?:;9I<  .?:;9n@�B   :;9I    :;9I  !4 :;9I  "  #4 :;9I  $.?:;9n@�B  %.?:;9nI@�B  &.?:;9nI@�B  '.?:;9n@�B   %U   :;9I  $ >  $ >  & I     :;9   :;9I8  	 :;9I8  
 I  ;   9:;  9 :;9�  : :;9   :;9  .?:;9nI<   I  .?:;9nI<  9:;9  :;9n  .?:;9I<     &   I  .?:;9I<  .?:;9<  .?:;9�<  . ?:;9I<  :;9  .?:;9n2<d   I4   .?:;9nI2<d  ! :;9I82  " :;9I82  #/ I  $ <  %.?n42<d  &  '.?n4<d  (I  )! I/  *.?n4<d  +.Gd@�B  , I4  - :;9I  .4 :;9I  /4 :;9I  0  1  2.G:;9d   3 I4  4.1nd@�B  5 1  6.Gd@�B  7.Gd   8.1nd@�B  9.?:;9n@�B  : :;9I  ;U  <.?:;9nI@�B  =.?:;9n@�B  >.?:;9nI@�B  ?.?:;9nI@�B   %  . @   %  $ >   :;9I  ;   9:;  9 :;9�  : :;9   :;9  	.?:;9nI<  
 I  .?:;9nI<  9:;9     :;9n   :;9I8   :;9I8  $ >  .?:;9I<   I     & I  &   I  .?:;9I<  .?:;9<  .?:;9�<  . ?:;9I<  .?:;9n@�B   :;9I   I  .?:;9nI@�B    :;9I  !.?:;9nI@�B   �   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  i_main.c    stdio.h   stddef.h   m_argv.h    <built-in>    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   doomtype.h    strings.h   inttypes.h   stdint.h   stdint.h   types.h   limits.h   syslimits.h   limits.h     	�@     ($sg[�vZ �   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  dummy.c    doomtype.h    strings.h   size_t.h   stddef.h   inttypes.h   stdint.h   stdint.h   types.h   limits.h   syslimits.h   limits.h     	]@     + {     �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  am_map.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    deh_main.h    z_zone.h    d_mode.h    doomdef.h    d_event.h    m_cheat.h    st_stuff.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    v_patch.h    d_items.h    p_pspr.h    d_ticcmd.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    w_file.h    w_wad.h    m_controls.h    v_video.h    d_loop.h    doomstat.h    dstrings.h    am_map.h    m_misc.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   doomfeatures.h    deh_str.h    sha1.h    doomkeys.h    string.h   posix_string.h   i_timer.h    r_local.h    r_data.h    net_defs.h    r_segs.h    i_system.h    d_englsh.h      	^@     �x;=/< .'  � > 
e..XY J&  �
u� L.&hc!Zd":	.g	�gY	�g	�e	.g	�/	;g	.i	/g	,g/eg&����&	"gg	rg	g0��tX<Xg-g<fhjce2
9egYsgXg4+�+t&< fu+'�&W fu"'<<h'�x�6txf
 rq�d��x( .ZJZ
�JL
�<.,	zfgeg	k7h	Y�/	� �Y;gZ,hCffh��	��	h	,hJf.
LfK� f.
LfK�g
fe
.g' vf
tuf��v<v�����Y	�g	�it	��	2�	0=. 7
ft�<fY	;g<	Xg[lTrghrg` z u  � � 9li$* P , 0 Y �]X# 2  � ;h�'#	��	�	�ZY�eg/��g	.#YW�Y�4# �Y� ��Y��Y_!gWgXg_!gWgXg
Xw	f�2 ��Y	W�
[�		>�-  �-  � X1�2  �.  �- X .��w	.  �-  � X1�r.  �.  �- X .����������XZ�ftg0YXZXZ���Xgt/����Xgt/���.�Z!v�� .�Y� � X � ��fX.<
��� .	L	>�f  J+ ���f  J+ ��) ������.J '#sgXhf�
Y�Z`�<" ��@ff$tX�fe$.�/sg$���eLdggt<
�^f�%�%tfg+ X9 �#f#<.�'�%h�[�[�]C�/tY e�<f
L�=W
L�	Kv.fK<
/�>JY<
/�>..@�<.Y��e=��=e�KY��e=���> J � t < . 
�* <   J� X t < . 
�* <   �$yt {zJjJ�wh	<;K	/	H&LJ/v
hK=	$=	:K$/<*<J/Z
v;K#	:#>	,>	;X./ /;=0
vK=	Kf	;'=J=22L=W= J � J < . 
X 
<2=W= J � J < . 
X+ <   �\Y�<& X tY< J tY<�<	��X�=c.&.tf@b<�NbJ @b< @9NE==Lfg�	g	L=0=x..f�g�	Y	L=0=.x<.  
X 	1XXKuY (z�g�u�-0	c�KfK  Z 	 V =	  K  j X2g�/u�-0	c�=fK  Z 	 V K	  K  j X1X .'$ .��b</�Hg/;gg< JZ+�	J^vvZ�Ih���K�
th	- X � <[  <p�..<Y�=�
a@YI=�vK ..<�8� N�/;KLLueKXMY"L:M8YKLLueKXMY "  � bJ < Y J L XZf....#yC�tYjy$. �# ���Ke1vH�. p�fPj* $�!Z*X<<1..#y�\�=	e��	 � <! �	 e! K% <? �2 �K� uJ�[fX.t<t.L#�#u��YY��Zv x   r  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_mode.h    doomdef.h    doomdata.h    d_ticcmd.h    d_loop.h    d_items.h    m_fixed.h    tables.h    d_think.h    info.h    p_pspr.h    p_mobj.h    d_player.h    doomstat.h    doomstat.c    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   string.h   posix_string.h   i_timer.h    net_defs.h    sha1.h     C    =   �       dstrings.h    dstrings.c    d_englsh.h     �   B  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  d_event.c    d_event.h    stdlib.h   alloca.h   feature.h   null.h   stddef.h   size_t.h   wchar_t.h   locale_t.h   posix_stdlib.h   doomtype.h    strings.h   inttypes.h   stdint.h   stdint.h   types.h   limits.h   syslimits.h   limits.h     	[&@     #t<<K-�!�g%h,�@!.b!N*xh �   �  �      /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  d_think.h    info.h    stddef.h   stdio.h   doomdef.h    d_items.h    d_items.c    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   doomtype.h    strings.h   inttypes.h   stdint.h   stdint.h   types.h   limits.h   syslimits.h   limits.h   i_timer.h    d_mode.h     �   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  d_iwad.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_mode.h    d_iwad.h    m_argv.h    m_config.h    w_file.h    w_wad.h    stdlib.h   string.h   strings.h   m_misc.h    posix_string.h   i_system.h    <built-in>    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   ctype.h   config.h    deh_str.h    doomfeatures.h    doomkeys.h    inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   d_ticcmd.h    d_event.h    z_zone.h      	�&@     �b@Y;u	\*v	W	< x� 	  J Y	  � � 0�{f	Z"	="-	�f�'z�x<	4X�\2�	4..J+�L�. .n.	]fZ:	>X	O�3.�
< ?Zv 
 
rtrX�JXZ	�t.	Z�	>Z�	[�}	�	:Z	ZMy	.f	��JuJ�X�	�\8ZZ"  �  �}�     �	�}.t	�Mt	�%J"�	L�4
�	L	�<?�Z	�O�	.Z>.sJ�<<	��B�Az^zXBz.'y.&�	.f	k	�Z <u -K tJ�?9�.<.'		0$J�t   <
fY#X	0) XZ.J$ ~ . J`Y#X	0
YZ.J# �$ U . J	XY �	   �  �      /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed /home/user/.local/share/lemon/sysroot/usr/include/abi-bits  d_loop.c    stddef.h   types.h   stdint.h   doomtype.h    d_event.h    stdio.h   d_ticcmd.h    sha1.h    net_defs.h    d_loop.h    i_video.h    m_argv.h    m_fixed.h    net_client.h    net_io.h    net_sdl.h    net_loop.h    i_system.h    i_timer.h    <built-in>    stdlib.h   alloca.h   feature.h   null.h   size_t.h   wchar_t.h   locale_t.h   posix_stdlib.h   string.h   posix_string.h   doomfeatures.h    strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   seek-whence.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   net_gui.h    net_query.h    net_server.h      	�*@     ��  	fzf
. � � <	 ,	f��{ #Zr0	3f�1 <�1j�Y��*�p	�pf<JOf" J]s.]]s=;K
<5�J?5+7�5�ut
.�k<Xu�hf	L�.u.	/
	z.	�	0XH.JJ 7�	Ze	ZXy"X^ X�	�3<f3 J3<5K3;5u3I5׺ w<f=u	 !"Xtg".� e�s=�	��#w	 wX	<XZ� <� � f�<v
�Ys{yt/k	0X2[�~%��~ft�% %<f2k�%.d<	<K./	]t?��~f�	��p<	�fZ	j -<g-s f	u�*�:�����0 38 � .�	Z�~��~ft�tY�Xt.	�o�XJ'.�Y � � � � =  j �~     � �~<	0s	u/&o.JX �  < fXXa.	�X	�!+f!X+t�r	v	�.	�	�	�	�	�	��+ �  �.<wu �   q  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  d_main.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    sha1.h    deh_main.h    d_mode.h    doomdef.h    doomdata.h    d_ticcmd.h    net_defs.h    d_loop.h    d_items.h    m_fixed.h    tables.h    d_think.h    info.h    p_pspr.h    p_mobj.h    r_defs.h    d_player.h    doomstat.h    dstrings.h    i_sound.h    sounds.h    z_zone.h    w_file.h    w_wad.h    s_sound.h    v_video.h    d_event.h    f_wipe.h    m_argv.h    m_config.h    m_controls.h    m_menu.h    p_saveg.h    i_system.h    i_video.h    g_game.h    hu_stuff.h    m_cheat.h    st_stuff.h    am_map.h    net_client.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    d_main.h    stdlib.h   string.h   d_iwad.h    w_main.h    m_misc.h    i_timer.h    i_joystick.h    p_setup.h    strings.h   i_endoom.h    wi_stuff.h    f_finale.h    <built-in>    ctype.h   seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   posix_string.h   config.h    inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   doomfeatures.h    deh_str.h    d_englsh.h    v_patch.h    net_dedicated.h    net_query.h    r_local.h    r_data.h    r_segs.h    statdump.h      	�/@     �g-�5u�  �� x� ( �O��t�x<�'�Z�L��.%t[.MZYYZYYYY�w�Y���������	   *	 2 Y  _X� .�m�(!K�}�q	�f��Y���-^��[%YjX��Yg-J"t�����g1Y1Y[���1p���#f�������\1��%���.�Yj	��lztg��"�i0uW1�
:�
Y4;:�<&Y\LXg<]0X>ZW;/�Y�	z<	4�YYYX� �! �7 �	���Z�Z�Y�YZYZZ	��ZZ��)t�((!&tqX%�(qfv�%�u<(���[&�#g�S���J�fZ��mXww
��1t�	Y��x� � K	�L�6���� ��  yC	 �Z L�		
o.XL�	
	v.�	��N��		.s�	�	Y�)t�.� X�X
	�	J�	J�$Ht\#f�2�	� � � �� � .� X� O!�W/Zd�	xL�~��f\�~��Z�~��L�~��	LL�~!���~!� �& L�~��Z�~��Z�~�� ) �  % � <	ZJZ��  x6xt�\��� X�xXn`xXn	XwX	fZ,h	X	�K
�	�K��	�t��
b\<Kt.X��	j�!'f!X'<<g!'�<g!�<g!�<f�[��Y[��x	Z����|t���xY�|
	�N.�	���XL.t�	.f\�\�(f\�Z�ZJ�f$X	��!X"��	Z��	�	L�>�=?8	Xs�f	Z
J�	�$.$XJt��x	��{�Y�Z�Z:0�	��	�?�X	X2px2�xt4/�L�K� H X	�	MY��R��z�	�/ J, �	L�[�YYY�`[	s����
�	ZL�X=��
	�L�X=���	
v�
�	ZLt.�
f	�L�	�	L�KX1'>*:>*dh0'X*<<�	��	�	L	�	�	��	�	L$t.�	���Z�Z�Z�؟ZZ�Z�^# �  �	K�	�	L��	�Lt.��	�L��1	�L�[f	L	XK����[	�y.�Z&JJZ$ �   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  d_mode.c    doomtype.h    d_mode.h    strings.h   size_t.h   stddef.h   inttypes.h   stdint.h   stdint.h   types.h   limits.h   syslimits.h   limits.h     	�C@     2	3) � � H�8]$	Z�.��.<JsX	<
KZ=e<Ju �& z� < Jf/%ih�<X	L<1K ?�	3
�� G	f8]%vt #�� �   z  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  d_net.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_mode.h    doomdef.h    d_main.h    m_argv.h    m_menu.h    d_ticcmd.h    i_video.h    g_game.h    doomdata.h    sha1.h    net_defs.h    d_loop.h    d_items.h    m_fixed.h    tables.h    d_think.h    info.h    p_pspr.h    p_mobj.h    d_player.h    doomstat.h    w_file.h    w_wad.h    deh_main.h    <built-in>    w_checksum.h    m_misc.h    stdlib.h   alloca.h   feature.h   null.h   size_t.h   wchar_t.h   locale_t.h   posix_stdlib.h   doomfeatures.h    seek-whence.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    d_event.h    i_system.h    deh_str.h      	�D@     � zjt�	� �. �v[O$But$JutOh$p�.�	0X Jnoy	/Z..I� XG6XGJ	xX�	X	L	�	�	�	L	�	�!kSK�!Y!f�xSO`!�?xXXJ	
XvX
f	X	L�_M	����fuXK������� ��Yf�� t�tJ� Y�~PzJgOgzJgOgzJgOgzJgOgzJgOag	L'�	J� .�tX	f�	f�	f� �f<f� w�f J	�  X � VQ!��� -   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  f_finale.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    deh_main.h    d_ticcmd.h    d_event.h    z_zone.h    v_patch.h    v_video.h    d_mode.h    w_file.h    w_wad.h    m_fixed.h    tables.h    d_think.h    doomdef.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_sound.h    sounds.h    s_sound.h    d_main.h    dstrings.h    d_loop.h    d_items.h    p_pspr.h    doomstat.h    i_video.h    r_state.h    hu_stuff.h    ctype.h   seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   doomfeatures.h    deh_str.h    sha1.h    i_system.h    i_swap.h    string.h   posix_string.h   i_timer.h    d_englsh.h    net_defs.h    r_data.h      	dH@     � 	
 \rX1����	��hy.9zu�"Y	v.% fZ	w � �
Y* J
gh K t pJ���� Jt.t�fY
r��t < = I �  ]  y����g'W<Vv� wZ	<YLZ	K1	1GX=^.�=<��
O4X0�:mw���:�M��y�z��`	��y't+f<�	��f��!'��Ku1u1�7J�u]� �5r��5;J���=e!6����%���6����Jut�xtowtq{^wf���J�9J�9J����0	HK����9?��	��W���}<$��� e��_�dhZp \�(�3JfZsd��/ZiX��.	-[	�i4s��4�:J�*xb!�Kr .�.�} �	[�<u6x<	X0Z	<gJ�.gr.X=Z=1.�=.6	<KLX=Z	=wX./s�KY<1  Dx(��i u S8/<8JX%tJK
#K>fZ�=KZX 	Q@     +=+�X=<L#�+gZt�K01	JX0'w
	.w�
	fY�=
Z
�>Z05f0�5X&�>���"7AX7�f�	v	�#�1 X�.i��iu�#f., ?[[Lf	Z\�jw	^x 	�J	k � =   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  f_wipe.c    stdio.h   stddef.h   types.h   stdint.h   z_zone.h    doomtype.h    i_video.h    v_video.h    m_random.h    string.h   feature.h   null.h   size_t.h   posix_string.h   seek-whence.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   v_patch.h    f_wipe.h      	JS@     � 9u80v<ZXJZ	0
/Jl0
/JK
h
K[<1>')<
v.

.vX	Jgt

X v. pt

 	<
rt>	<	Xg�\<� >Z	JLfZ� � =  < J  ./ (; g(I�+<Y& � v  � K Z#/ =:K!<Y &J�. f Z  � K Z.<yJ�~t+>,t�� !tY���~J#�.#X<.XZ �� � Y  � J X <Z�0> ..,X 	�U@     � +*+28@xx. 2x\��0xf\.uX�� vY
�
!�=JJK J �
V L  f1J� <!.XXY;uYRY-=W=WJKY;uYgt .
 w.	��u<U�u��<L<����=... n!   .  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  g_game.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_mode.h    doomdef.h    doomdata.h    d_ticcmd.h    d_loop.h    d_items.h    m_fixed.h    tables.h    d_think.h    info.h    p_pspr.h    p_mobj.h    r_defs.h    d_player.h    doomstat.h    deh_main.h    z_zone.h    d_event.h    m_argv.h    m_controls.h    m_menu.h    i_video.h    p_saveg.h    d_main.h    hu_stuff.h    m_cheat.h    st_stuff.h    am_map.h    v_video.h    w_file.h    w_wad.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    i_sound.h    sounds.h    s_sound.h    dstrings.h    r_sky.h    g_game.h    i_timer.h    i_system.h    m_misc.h    stdlib.h   m_random.h    r_data.h    f_finale.h    statdump.h    wi_stuff.h    p_tick.h    p_setup.h    string.h   feature.h   null.h   size_t.h   posix_string.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   math.h   seek-whence.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   doomkeys.h    net_defs.h    sha1.h    doomfeatures.h    deh_str.h    deh_misc.h    v_patch.h    r_local.h    r_segs.h    d_englsh.h      	�W@     �X?�  w$JUw<.qf$�9>I?u5�&t � t�
w�
tY ��u��%*	��	Y]Zl.M<vM<vK<�./<t3K!<�K!<�KUt+.K.T,X/tMPt0<��t�
<�	�<�.	/<�t�t�t�	�<wt�t�t�	�<�X>t. � t�t�Lt�t�t�L
�. � �	��~�	ZC3.	O<�:,^�yJ:x�+<.&t:B�+<t#	.K...J<=X�t#XQ<Y<5,t�K�f(	�=sX	.�<�<"=<Y.<	 xfq�tL
<�t	��	�8 �ZgKg�K���Z�	�u � t	�% �ZgKg�K���Z��vfYJ0�	N!��d�.
Z�
Lw/?��M��:f+<k	�,	�-4f#3)	O#t.X.Cw	 �pj$/�	�V\	Xfhrh/��V2s� .g u En�g�g\�[)zt�/�W/~����#���0	0(�=.� JY �- J9�a/	Y/<(  	�� X� Xp"  ��. J��Y]Jx��������� �	_#4X% J  J	�
 �% 	�
�?����Ju	�w�Jj5v	f5<Xx�	NZN�0D�<nf�� &)f&X<)f	<g)f	<g	[�~J
x,t	f,3X	j�N\�0	D<t<l�<g	��	_.�.t=s/�t���	 B�quv9v0u 'zsfv!u�vx��y�����h� X 	�c@     � y5y�_t w�$�(<	< Y$J<
Yt<2=s
9=>
JXNfY�
�:Ft&<!�
HX
fX	<Hf�	>2gg.
�ggv.gg0gg	. t<=u0�.	1.J<!X<����Y	���J=YXzt
fY-KXL*/*;K z. <.�X-_��st�pt  #0h�\f<�	J
J	L#</=:#JuYy �<Xs<f>r^� ��$�#��/�-J$#��� :j�Z�	\�|�uX�� �.`�����.f��<iZK�#�W#�2?4K�
[����y.�0�5i����Y <
�Y,t	�!�|v�h Z  y s � /  @ F =  g  g  yf�U��ZY`�	fK#v��	�\#"e�.gY��. =�Y�=."WgXY�1zO/Ye=^z�BXv	\"�"�	=X	uZ���YYYZ]# �  �	���	](����Z$x  $*#Xggg� ��	�!X�	�	m	N^qtX. TXMZ�*^ZW f�� �, f w  f I�!��
 �$  w  f I�!�� �  pt yf �  �  �  �  �  �  �  �  �   g  v  	0WZ	2x< Xi<I�}X%��Xv��
X	Lt	e \iZiYYYZ
XK���[X� .
 w ����'������Y��.&zf_,�.fK��utY
	�Kt.
�g��;uvNkأw�$�	X?w	 )�tjfh�	0�	\X 1 � � � � � � � � 1	  t	 � � -h
.u�* 4z�3�ZHvt>X	L
�	[	�
� V	^"	V0$t!I=uIKu	IYt��������� 1    � ;i�
�
 � �K�Qs�Y�\ �h-�&y CX]vy h��� #	�	YemU+�I	/,�z J�PJX	��
vt�
�
��$�����	�/v	Zw	fL	 =,�,t<Y���[/�|.	t[[-�K*�jJ!vr	0#KI	K#t'J<	�5J<M* .=# qMw/ZvJ�/tX�2	Z�	/t	�J�1X�rvJ	Z�JsJ`��rL<s<*Y�a=*<@2�u;ut1=<IX 	�v@     �wz�# � t�t :kh:L�Y0Y0Y0Y0Y0Y0Y0Y0�,u,�!6	f�	t>>�t	�r	v/�	�
�h"�fK!<�K��0"u0�!	 �* � �L�$<J�Z�JY>J< Ot9��t	fL�
�-g
/vx
�@+u+�� f<"�) �	�[�.X+qXYYYXq.\Xu.\Xy._X :
   *  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  hu_lib.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    doomdef.h    v_patch.h    v_video.h    m_fixed.h    d_think.h    tables.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    hu_lib.h    d_items.h    p_pspr.h    d_ticcmd.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    ctype.h   seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    d_mode.h    doomkeys.h    i_swap.h    r_local.h    r_data.h    net_defs.h    sha1.h    r_segs.h      	�y@     $#YK�	 s
X/r
J=
KKmKJ&
	K-\g-YY	Wu#<.M	0V�u&x	Jw<|/w 	<h�u=�
fuK	<�Y;Y2=	�<4	YJ.vZ  ..,Z  ..Aw	��
< �'  Z m.�hK;=sX=,  fL	f. J fK��f&Jf3yX=.t..f
Wg:�u�  Y  ; u
 �~J >' �J �~. �J �~J �J �~< v �t �~<  
  K   m     .�#	f	f.���~�uKt� . K  t �0'�Y	YJY4t<�JY-t<�#
tb � fL�/
 0   ? w. 4 J ? X1. #$* \� � tY � t �0�h. 
 �~�XK�~
J�.��~
=
KKmK�Jx%�Y#=�<u$�~YK�J�~t�J&gJY'<<ug( 
=JZ<Y�0K�q	XA #
JZ�#!s= . JYu<Yfg  �	   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  hu_stuff.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_mode.h    doomdef.h    z_zone.h    deh_main.h    i_video.h    d_event.h    hu_stuff.h    m_fixed.h    d_think.h    tables.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    v_patch.h    hu_lib.h    m_controls.h    w_file.h    w_wad.h    i_sound.h    sounds.h    s_sound.h    d_ticcmd.h    d_loop.h    d_items.h    p_pspr.h    doomstat.h    dstrings.h    m_misc.h    ctype.h   seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    doomkeys.h    doomfeatures.h    deh_str.h    sha1.h    i_swap.h    net_defs.h    d_englsh.h      	�~@     �x 
t  �  � � 9li�#A�t�{y�{zX�����^sgIy �.z�z�.�0���		���<Y'X<ws�YIz  �[�M"���vZ1"��Z]	zf� J .����
� Yʻu��� g �g�	�	/t�g�t/
�)�f)t/��
u"T���
1��� _<&�
��<�2uh#my.�=.;gn#p<<
�.v
tg[�����0
 � <��XYXVZ Z c t�ffk��
 ����<�L/Y	�Y	�Y	�Y�� i<W<� t�=	M?U�W<Y!</����Y!\>X�/	M�	hs�0="?g� k   e  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  stdio.h   stddef.h   types.h   stdint.h   doomtype.h    i_sound.h    sounds.h    m_fixed.h    d_think.h    info.h    tables.h    p_mobj.h    info.c    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   stdlib.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   doomdata.h    doomdef.h    string.h   posix_string.h   i_timer.h    d_mode.h     �   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  i_cdmus.c    stdio.h   stddef.h   i_cdmus.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   doomtype.h    strings.h   inttypes.h   stdint.h   stdint.h   types.h   limits.h   syslimits.h   limits.h     	        &/B#!�� �   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  i_endoom.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    i_video.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   config.h    strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h     	p�@     $+ �   5  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  i_joystick.c    stdio.h   stddef.h   m_config.h    m_misc.h    stdlib.h   alloca.h   feature.h   null.h   size_t.h   wchar_t.h   locale_t.h   posix_stdlib.h   seek-whence.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   doomtype.h    strings.h   inttypes.h   stdint.h   stdint.h   types.h   limits.h   syslimits.h   limits.h   d_event.h    i_joystick.h    i_system.h    d_ticcmd.h      	r�@     � 4�.#� t.MY�������	  * �	 1 Y � ^X �     �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  i_scale.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    i_video.h    m_argv.h    z_zone.h    <built-in>    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   stdlib.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h     	        � s*u;K<*o<=
;u*7<=.Ju>JXc  	 < J L  J J!  Y  J J"  Y  <	 0 s .	 = 	 =  t qJX  s*uz<AKz&<*l<=
;u*7<=XXuK> P	 h �  ? 9 J! ) X1 / J Y  J$ " J) X0  Y  J J" ) X2 0 J Y  J	 0 	 = 	 = 	 =  t n .� X <s*uz<A�z&<*i<=
;u*7J=<tuKK>  �	 	. J Z  J J! ) X1 / J7 X=  Y  J J" ) X2 0 J7 X>  Y  J J" ) X2 0 J7 X>  Y  J J" ) X2 0 J7 X>  Y  <	 0 	 = 	 = 	 = 	 =  t k .X f<gz4zt*5y<*5yJ4z<75=<yJ*P==<*s>9
=uKXYX�,;YZ J ��	 Z   A 7 J! ) X1 / J7 X= E XM K J Y  J$ " J) X0 7 X@ > JE XL  Y  J J" ) X2 0 J7 X> E XN L J Y  X$ " J) X0 7 X@ > JE XL  Y  J J" ) X2 0 J7 X> E XN L J Y  J	 Z       t h .  f.J�<	 A - X% X+ < X <	 K    7�> 	 3  <	 = 	 K   7�$	 4 + X# X) J f	 K 	 K 	 Y    y<	��  	 3  ? G	 = 	 =  f	 =  z�$	 B + X �# F) < X	 = 	 = 	 = 	 =   x
��  	 3  <	 = 	 K  <	 K 	 K   y<	�$	 4 + X# X) J f	 K 	 K 	 Y 	 Y 	 Y    w<�� 	 v  3	 K z<	 = 	 =  <	 = 	 =  <	 =  x
X�y )	o2*y<Cyf	<)8s*.
<u)6<<v 	 Z �	 ; /   b <5X� y5y.�yXQyXQA`xXh�A^q� f   
 S< =" ,f+ f: <( X < u " J+ f: J( X < u " J+ f: J( X < Tf ,. K H        	JYW=WK=IYXeKI<	?<2�u<.J�!-<J	y<� ��� J�X,.1 f{s6.tr*�u	w!	#��	?�9 <	��9	?t� <	�	?�9	?�9 <	�f9	?� J	�	?� <P4�L 4XA�?<, ,.1 f{s6.tr*�u	w!	#�	?��	?! <	�	?�	?��	?�9 <	�	?�fq	?� <	�	?�	?�c	?�9 J	�	?�	?�t <�� �� � X��� <. ,.1 f{s6.tr*�u	w!	#�	?�	?��	?� <	�	?�	?�	?��9	?t! <	�	?�	?�	?�9	?�9 <	�	?�	?�	?�c	?�9 J	�	?�	?�	?� <�� �� � X��� <� ,.1 fy
uvr!j x$t�nd<	z(7Jt,qJ2<$X<	@(7J,J2<$XJ	@(7J,J2<$XJ	@(7J,J2<$X<	>kX	.	=�	q.<�  ,.1 fy
uvrW.
ttJ.� 	V�L4L<	z	=J&J	ZJJJ	"1J&X,<f	KJJ		KJJ	"1J&X,<f	KJJ	"1J&X,<f	KJJ		KJJ	"1J&X,<f	KJJ		K�	S�	� 	=	�w X	qJ<< ,.1 fy
uvrfJtV *tW�;XEJ;<	:AYL'	_X	>	oJJJKXX\#2J'X-<f	LXX\	LXXYXXZgJ�	9s	=	�w 	Xqf<�  ,.1 fy
uvr�f�� V.*t� =X5t �JW=� <	��YK� �t	z	=JJJ2J	NJJJJJ	JJJJ	JJJJ	"1X&X,Jf	YJJJJ		KJJJJ	JJJJ	"1X&X,Jf	KJJJJ		KJJJJ	JJJJ	"1X&X,Jf	KJJJJ		KJJJJ	JJJJ	"1X&X,Jf	YJJJJ		KJJJJ	JJJJ	�	G�	� 	=	�w X	q�<* ,.1 fy
uvrhJtk��X WXY;>'<	:RYKktL		=JJJJ=XXXXKXXXXKXXXXJv<�	%s	=	�w 	Xq�<�x ,.1 f{s6.rt*tum	��	s/�	MK� <	�9 <	�� <	�U J	=	;/ h�d X .Yt'<�~ � XXY��Wut��YuX&�&XXY��YuX� ,.1 f{s* u6y	w�	w9	?�	?�	?�	?�	?�%t <hX	�JW6X	u.,#l,zf#B,z<#Bz<	v.�:0	<JS6<�x uug�  =t	ZY����	uXwt	ZZ��v  �     �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  i_sound.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    i_sound.h    i_video.h    m_argv.h    m_config.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   stdlib.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   config.h    doomfeatures.h    strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h     	,�@     �w	.wX	.`xXD`xX6\ X	�L
e�	[L��	� L��� 	v.
J <#t	Z	#?t	ZLTt	Zyt	ZB?t	Z	#?t- X J	ZTt-XJ	Z<t	Zi	�	�tX>#t	Z`	�	��fB?t	Z>#t	ZB?t- X JZ0#6t	Z>#t	Z>#t	Z>#t	ZB?t	Z>#t	Z>#t	Z>#t	ZB 1   �  �      /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  i_system.c    stddef.h   stdarg.h   <built-in>    stdio.h   types.h   unistd.h   stdint.h   doomtype.h    m_argv.h    m_config.h    i_sound.h    i_video.h    i_system.h    w_file.h    w_wad.h    strings.h   m_misc.h    stdlib.h   string.h   alloca.h   feature.h   null.h   size_t.h   wchar_t.h   locale_t.h   posix_stdlib.h   seek-whence.h   ssize_t.h   posix_stdio.h   off_t.h   posix_string.h   uid_t.h   gid_t.h   pid_t.h   config.h    deh_str.h    doomfeatures.h    inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_joystick.h    i_timer.h    d_ticcmd.h    d_event.h    d_mode.h    z_zone.h      	e�@     � MUMZr==Ku. %�  0h8"V >.$�<0 	 Y W	 = X0=.-\ 	 ] � .3Y\JYY�Z�I
.<%v	Z/J6 �  |	��{���	�wXLY��:�V�K��Yv	Zh	?J1��~�	��~F�8�I��8=LJ	
J�ZY	?	K"o	<<2x1IK��=�[��� �  �}.u	.uX	JuX	fZ	L"t.�	/A	$X	>	�Z	pr<��[X.� [	�XtX	�X	>�#.#�<#J��L��L��L�D>. �% � ] � Y,  v�f��X	r.2$�	=03<u4<AJ3W%K	g01:u=2;K?I=#<1,#h:/2<?J#<	Y\X 	 s   �  �      /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  i_timer.c    types.h   stdint.h   doomgeneric.h    i_timer.h    doomtype.h    strings.h   size_t.h   stddef.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   stdarg.h     	}�@     %	xw	t		�hht</6d	i t	�hg3X 	Ӎ@     $ \   H  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix  memio.c    stdio.h   stddef.h   memio.h    z_zone.h    <built-in>    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   stdlib.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   string.h   posix_string.h     	        *	Mq	MU	#Z=K�. %h%XY
J.$rf,J<:<$t<Z	<]<<<jJL%	#�	�>Y�=�J%
OEMnJ�>)J!<fZ��=/�=f<�<>gM�<=
J=#!I=0<[=X 	        =#�yJ=1=.h=
5e Xu
> �   *  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  m_argv.c    stdio.h   stddef.h   doomtype.h    m_argv.h    string.h   strings.h   ctype.h   seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   stdlib.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   posix_string.h   inttypes.h   stdint.h   stdint.h   types.h   limits.h   syslimits.h   limits.h   i_system.h    d_ticcmd.h    d_event.h    m_misc.h      	Ս@     +yo?c#X. <L�Xj=� J 	$�@     z!Y�� %q#�	^L< E   �   �      /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed /home/user/.local/share/lemon/sysroot/usr/include  m_bbox.c    m_fixed.h    m_bbox.h    limits.h   syslimits.h   limits.h     	[�@     #��'Y
YY=Y
KK/ �     �      /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  m_cheat.c    m_cheat.h    stddef.h   doomtype.h    string.h   feature.h   null.h   size_t.h   posix_string.h   strings.h   inttypes.h   stdint.h   stdint.h   types.h   limits.h   syslimits.h   limits.h     	��@     %b@ff" Xg>J	^+g	�
�<	]3	>3,	Z?<g	h1vV	�&=�</ (   z  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  m_config.c    stdio.h   stddef.h   errno.h   doomtype.h    m_argv.h    posix_string.h   m_misc.h    stdlib.h   i_system.h    string.h   seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   ctype.h   errno.h   config.h    strings.h   inttypes.h   stdint.h   stdint.h   types.h   limits.h   syslimits.h   limits.h   doomkeys.h    doomfeatures.h    d_ticcmd.h    d_event.h    z_zone.h      	8�@     ��+# J	Z/</f��l/tJ� %7AS3X>	Z�A	Z�[X �~ M X	g	J��v� �uu'�~��~�'k�~��~�'s	 �L!�!WY-u	x Xw	.	�	L)	�)W	Y!-	u	u ] Xw�� ��  . ?ZKu &iX>,& X <O�}�J�~X�)J'�=2'J%�/5�y.=Z.{%&I=%/11'�)J��Y<%#Z+ XgkJ/M#Z+ XgkJ=[#Z9 XgkJK.#	Z	�fXY[w	t	Z�u	X
tZ	�b 	��J C   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  m_controls.c    stdio.h   stddef.h   m_config.h    m_misc.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   doomtype.h    strings.h   inttypes.h   stdint.h   stdint.h   types.h   limits.h   syslimits.h   limits.h   doomkeys.h      	p�@     �!���������������������������\!���������\!�����������\ w�������Y���������������\!��������������\!������������\!�������������������������\$T2T&z.NZ 	 Z g � X0X ( �   k  �      /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  m_fixed.c    types.h   stdint.h   m_fixed.h    stdlib.h   alloca.h   feature.h   null.h   stddef.h   size_t.h   wchar_t.h   locale_t.h   posix_stdlib.h   doomtype.h    strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_system.h    d_ticcmd.h    d_event.h      	��@     $<<(Ju	 
.
.<
<fJ<.LJ�<<	LX    �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  m_menu.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_mode.h    doomdef.h    dstrings.h    d_main.h    deh_main.h    d_ticcmd.h    d_event.h    i_video.h    v_patch.h    v_video.h    w_file.h    w_wad.h    z_zone.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    hu_stuff.h    g_game.h    m_argv.h    m_controls.h    p_saveg.h    i_sound.h    sounds.h    s_sound.h    d_loop.h    doomstat.h    m_menu.h    m_misc.h    i_system.h    i_timer.h    ctype.h   string.h   <built-in>    stdlib.h   alloca.h   feature.h   null.h   size_t.h   wchar_t.h   locale_t.h   posix_stdlib.h   seek-whence.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   doomkeys.h    d_englsh.h    doomfeatures.h    deh_str.h    sha1.h    i_swap.h    r_local.h    r_data.h    net_defs.h    r_segs.h      	�@     ��ht/!>!"��~ &��XK� �"���!�!���!���}�wX���t�8�AW/g9�/J/Xt�
�Ku<g� JDb��1Gt	X9XYE;XF.	X+XUt	X4X	X��uu. & �MKMY�$�MKMY�� $d�hZ�!>!!4�MfL/-g2fZ/-glJf?fKJfY�D ������Y�<�|X�#fYvX� �$����w�.�  ����x�K��xX�{ 	'	t�	�Z! �0K��< sJ�� \T 2W<uW�   � L : � _�L> ,X 	��@     <J%=J%.tY��t�t�t�/g + �#fYvX� �y<]SkS3XY;=;Y  Z  � > X g I �  .v�Xf�	��.<..,X 	��@     �| !�"%�t�%�tv,�� !�#	5�!tt5�!tt�*�t�)�tv,��LV>V4!=)WJLv>`LV>V4!=)WJLv>
Xhs�gug��{ ��tL�;tJ ;tY����tX��� <i
`x [U	�wXM�ztB���~�Z�Xy'/��w��.��(3a", A. �Z�=Y<0.�<.<1< DwzJ?LI/�. <Yu$ , <3 x	.w<	�v< 	<gLZ	=	<]	[G=^.�=<��0....�y $�#+$W# (  t �  t q]<J#�#+#�! (  t �  t q^�#0�#;tY#tXvL,X�
J��e�u, w�q�hs4E5X�����< � <ZJ��h#[K= o. <.<��M0�Y0s=0;.K;uYt���YMx*	>:u� 	L"hN� Z  � <3	1�Att1tAJ<���	 ;uu�t ��Xy'XY9X��X�v
 XYX ���v
 tLYY��,;J;tY���rt�	0
YQzt<. ��Y_	] �* ��f���}���. �! X�
Ld3	w
	X0
gX�h
g0
0
gX�h
gX�h
gX	�[f%.< � X�gX�* � X�e�;g	LgX��	K<5<LgX��
fie�;g	LgX��<LgX��
fi	hgX�	<ZgX��� J	�=A��M	f�,s�,3)t��)�Z[#s�#<	J���X>; �   s�t�$��*.<K*,g����) ����t�.0] �+ �K�Y\��".2�"XY[�Z�2�Y.�uZ�Y.�uZ�Y��[�.Y[�tYYZ�.�uZ�.Y[�tYY`���/%iqi'%.'tX�]�YS	� t
u -*<	.L=� Y(��
��
v	:Y!tL� Y(��
��f- ��.�$�t$.
��f- ��.��$X�
���t<$�J$ �- -�K	hu�/
��!��~�
��t�J�u�
	t�|J�f��#t	t#< �Z#	�/ V . . ..
uXu
p#	. r��wXX>X ���X  � w  U/Z$X!fKLX�t��Z1	gY XX=X�l�% �	 w% U		.X�X	����'�d�ud��
<vtg����2sv�w���x       �      /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/sysroot/usr/include/sys /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/ansi /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  m_misc.c    stddef.h   stdarg.h   <built-in>    stdio.h   errno.h   types.h   stdint.h   doomtype.h    i_video.h    v_video.h    w_file.h    w_wad.h    z_zone.h    stdlib.h   i_system.h    string.h   posix_string.h   strings.h   ctype.h   stat.h   seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   posix_stdio.h   off_t.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   errno.h   stat.h   stat.h   uid_t.h   gid_t.h   mode_t.h   dev_t.h   ino_t.h   blksize_t.h   blkcnt_t.h   nlink_t.h   time_t.h   timespec.h   types.h   id_t.h   pid_t.h   suseconds_t.h   fsblkcnt_t.h   fsfilcnt_t.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   deh_str.h    doomfeatures.h    i_swap.h    d_ticcmd.h    d_event.h    m_misc.h    v_patch.h    d_mode.h      	��@     7� 	ȳ@     #�	Z�	{��5JA[�?Y�?ZJ .'\TNX>.[/;=Z�  DyS�X=Y�]��>Y�=Y;=ZY�=X.... !WKWK	[�	 K	  K	   � .  #3a�.<	<[]� qJh<.XwtJ	�h�y 5 y._  . K  <	 Z   V > <0 	 z4zf�u<BY;uX�y	0>	.#�<� H <S<�iX>	Z�.@f�  %J	<	Y_	yJCtgY<< �<1.l<wG19M9XR737uXg		�	]I	K+�<y<.�=<	ZtY6	�X��;Y =y<<f=<<<2
L�.Xc?.uy<<X 	*�@     e=X<tX	� V L Y	  �<%e=X<tX	g V! " < �	  �<&z4z.��zJ^z<�0	�u.h		-	]�zX6�	ZtY1��		*	]z�.� �}<m<�t 	�@     �,UJuf\J<	Z	Y<.  $Q�W�Y }    !   �       m_random.c      	��@     2�<gu#�<gu#�� �   S  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_ceilng.c    stdio.h   stddef.h   types.h   stdint.h   z_zone.h    doomtype.h    d_mode.h    doomdef.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    d_ticcmd.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    i_sound.h    sounds.h    s_sound.h    d_loop.h    doomstat.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    r_local.h    r_data.h    v_patch.h    net_defs.h    sha1.h    r_segs.h      	�@     �3�.�  7n( .A�-J�Y�. y<
f�~.i{ y�kJXJZ��� � � < � S<	fJXJ[uX��jJXJ\Z�]JXJZvu.	.0Au	.�.3�(YJYh#>#�= y<f�~ v<
] X q� yf ��tux=�K!�Kv�g/>/HYs=2;u?!=?q�2�s=uKK:=X(X�< <..� <	21�(YJY<L&=
.V�#u w<f a
   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_doors.c    stdio.h   stddef.h   types.h   stdint.h   z_zone.h    doomtype.h    d_mode.h    doomdef.h    deh_main.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    d_ticcmd.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    i_sound.h    sounds.h    s_sound.h    d_loop.h    doomstat.h    dstrings.h    <built-in>    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    doomfeatures.h    deh_str.h    sha1.h    r_local.h    r_data.h    v_patch.h    net_defs.h    r_segs.h    d_englsh.h      	)�@     9�*�MuJXjuJXJ\uJXf��uuX
H$Z�xK;�YJX
fuu^
.h�uJX$J dX�Z��;u=3K;�	w 	X  �  x!._��E	4z.(��tuy	=�L�KKuv���IKU���Is�j=uH=yu�s�	YJXku��	YJXJNXX:X< <..�~<v�Jx 2 fh�5 fh�5 fi�X.YIY.�  Hv ��" fh�5�$ fi�5�! fh�tPX7XI7.	X�JZ{	g��+J�	� ��^%�J�	��;=YK�!zf�K�(uo�u4u�1uu��  . 'Mq#U#��Kh!�Ku�u. 	 Mq#U#Z:>ZyXK;zJh!I�uKY��.  E   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_enemy.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_ticcmd.h    d_mode.h    doomdef.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    i_sound.h    sounds.h    s_sound.h    g_game.h    d_loop.h    doomstat.h    m_random.h    i_system.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   stdlib.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   d_event.h    string.h   posix_string.h   i_timer.h    r_local.h    r_data.h    v_patch.h    net_defs.h    sha1.h    r_segs.h      	��@     �	W��ti:�
��Y<��[m �HuY�2<@ �w �Yy�.r<�t =r=Lh����f!t�Y#f��	Wj.X<.. J  Ig,u<X 	N�@     
@t	YJ>��0t�M�Pi�	KvfN�	��sue
cl
dZZ�Z�\y�;ZZ[�"��+]	X� 	< uJf	Yt>Y�"w"9=0)t
�);
�?Z,0fif�	<i	c/j�Wg1��yf�L	
2!f.4zXjFj/ht 
=XO"X�Z &u�Xvir�8K<g>
vu�B�
�c�n$0.$.0f(f.�g, X) �t�
�X	Xu.<<<..t���hu��
fx�v��L:hX�	XoXLPh�z�,\	th�zJ,\	
tm�u��fh�c�i� �X<.Xx&JZf��
/ v   ��Bt��MtXt�	ot	��
s�1_<4���".X<.	X�t�x t���7 x� J.hJ�uYX $F?�
vX
�r��v��sf
	Xf
�#X�=z.#X�=lz<;\1X't=� 	 #c?K�	�LY���fZ)=;YLKu	�Y���$t]fL/sg  f�8<H ]tg�L�K�$t<-<S ]th� ���M$t��^	�x���L�l�L�tgXZ�� 'tW\&:v�XAt�tX).<<..'��x(YK��>YtX/X%W?,==/Y .,/�$y�
.[sffnf
Xv
 Y�K0    t X /+ W > e  =   = - / � <4. J.. #z�	.wX	tw	 Y�K0X#."X/X.W?,==/Y .,/�$ >Z	X[t\$t>��N $ >Z	X[t\$t>��N #�N[��(�PY	�L�YY�<	.=Cy ^�X%�PY	�LYY�	<u>Z  #�PY	�LYY�<	.=Bz ]�X$�NY��%�P	XL�YY�<	.=Bz ]�X(�PYu
=vgg�  %y�t�Z
�
p@X�<K�
v ��<L��I�/I�BKsK/�=��?[z
z<L<X"f<t??  <$�MY�X$�PzPZ	�LY�KY��F<	.>>ZX 4 t�t�#t
	twt#<<#>�9hihduuucKKK> � <���su;uYv�tv�;ug:Kg�. .... a  < V < X=.�X 	7�@     � 	A�@     
yu�t[
�ML�tJUL��=I=Z:=;K=. .-Y<^X!W=Y=X 	��@     !W=Y=X 		�@     #�PZr$u:u�X
 ��y'Z
���g.(t
\(p< (t<>TD"Jx�DC"/;� �= sY"JY ��.<-Y.f  =Y�X 	_�@     k[u��=�
/<hr==5/;!s=�=. #kZu��=�
/<hr==5/;!s=�=. #�Z
��>
X=<hr==5/;!s=
��>
�<hr==5/;!s=�=. ..
 Ot�����=�=��=Y�=YW
r�2)t.X:<<=Xu1���/J3g�".7f^Xt<b" p>H<7<:j�<Y�W=YZ9Kh
��?
XM�  ..z.\�;u  ..-X	 �NYgX%=�":� <tA�g� 	g�@     	#q?t"X�=z."X�=lz<;\2Y $� 	��@     �KY%x' 	��@     =�Z�	f	��� t�f	0	�"Xt�%��%�%��&W\ �F�.� # � t � ;x t���7 x� J.O1JZZ	f_	Zu{f�z�u�Y5�uY 5 YX$!W=Y=X 	��@     !W=Y=X 	��@     !W=Y=X 	��@     <X_<XXKWY<Yg X 	&�@     
�uG� ���$=$-�v.J.�tX 	��@     t]z�qX4$ � �L�Y�<gX=Z��ZX�<g>w<	f�Y/W^zzJX .Y;0,V
?q=<
gt=Z�hZX�<K�  @X 	��@     
�
sgyfXu 
��#&.#&9fi�*s=<4<t$JLUi.X y�
Jv
.t[�?��	\W
ZW
ZW
ZW
vW
vW
vW
vW
vW
v�	��=	XK(t��= XF !W=Y=X 	h�@     >
rZ3�X  �
   R  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_floor.c    stdio.h   stddef.h   types.h   stdint.h   z_zone.h    doomtype.h    d_mode.h    doomdef.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    d_ticcmd.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    i_sound.h    sounds.h    s_sound.h    d_loop.h    doomstat.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    r_local.h    r_data.h    v_patch.h    net_defs.h    sha1.h    r_segs.h      	��@     0f�|�x<	XJ/
.Y.�<	<L/
�.h=6/
u.h
Z=
.�N J	XJ=
.Z.0
ZK�{ J	<L=
�.0K
�x=
t/  C#9[y�JXJZZL:�Z	f
LJ1uy�J[.JX. 	 w#	R-v���wU?2
=�K�K����9K���9K���9K�WL	����9K�Y&K��[�K�3�K��:G�K�:x:G�K�:XL[:G�K:W�L'�&=IYY\�l,K� h	�	L	�XY		�XY) t .. J;M[�?z.K�WL� h�L
�&V
�X
�Jh��' i. .�~.��J.  .tm.q<	.n<tr< o<XJ��twx
=�K��K_Ȑ*gm	?FK	=LjfBzt .�����Kw
>y.�Z:>ZpXXk�<Ko <�umJKKKi<X<XJ<..... �   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_inter.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_mode.h    doomdef.h    dstrings.h    i_sound.h    sounds.h    deh_main.h    doomdata.h    d_ticcmd.h    d_loop.h    d_items.h    m_fixed.h    tables.h    d_think.h    info.h    p_pspr.h    p_mobj.h    r_defs.h    d_player.h    doomstat.h    m_cheat.h    am_map.h    i_video.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    s_sound.h    m_random.h    i_system.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    d_englsh.h    doomfeatures.h    deh_str.h    sha1.h    deh_misc.h    net_defs.h    d_event.h    r_local.h    r_data.h    v_patch.h    r_segs.h    p_inter.h      	�@     � ��YXvf/ff	E|tYJ0��20�	W�w	xJ`0	���	nJX1	��	eJX1	��	\J$X0	��  	�<� . � �$ f�JtY�Ju��M�rv�Y��u.\KX0X�L,��ZwXKXX 	=-[/[9�hY 
=	-[=V> .Ji�u
 Lu1Z;u�1Zu1Zu1ZXYu.	=eiuY hCk�.Xx<|2��� ���� [��� ���� \��9?g�[��EA/u�[��9?g�[�;uX9�Y�]g�.<Y���~Xg�X4g�X4g�X4g�X4g�X_X<X��[X<X�g���~u��[�~X<��~XY��~Ju��g��~;u���1�~u��1�~�u��1�~u��Y\yX�J<	X��[.�X��[�<X��[�<X��[�<X��[�<X��[�<X��[�<X��[ �  t Iht 1 � / WZ�\t<X��[�<���[t<X��[t<X��1t<X��1�<���1�<�L�Y1X�}t�X�g�su�YK -YJ 
 $b@�rh/�gIw9gt . t[gh�*3�
h �ji[Y*3�L>:�uZ<��]!tX�<O�X�<h	<wt	f6�xx_
��  fy�
�v
J��0-�wu ��	4��YtY�f�J0]oA	fwY��JuXL
uMsK�=�@�J<ufLB���XL	/W1	�	XM�/-Y�~]S\��<Y?�?��LeJf  ..eJ\XtYfh>dh[r� .���%ru���<KG?  ..G�X� �X� _   !  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_lights.c    stdio.h   stddef.h   types.h   stdint.h   z_zone.h    doomtype.h    doomdef.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    d_ticcmd.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    m_random.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   string.h   posix_string.h   i_timer.h    d_mode.h    r_local.h    r_data.h    v_patch.h    net_defs.h    sha1.h    r_segs.h      	0�@     �[+J<JLu\K<<� �J� ZK�J� ZKx�} UPZHZ3J:>#.M.�u  & [+J8NJLuX\KX,<[  S Qyt3hXZ:>ZIL"9�=YKsg. ( Pzt2hXZ:>ZIM"8�>X=�X/<Y. * [U[+MU1Z:>ZFK8Ku"�=X>YwhYX<vu. ..'\8%�Ltuw�0   (x
tv<Rv ��
K <h
K�ZJX<1! rJ+ < J. X.
 y	tw<mv ��	 vhK�
[JX<2 kJ& < J.  J.# 	Mq	#U	#��K�=K�=vg.  �   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_map.c    stdio.h   stddef.h   m_fixed.h    types.h   stdint.h   m_bbox.h    doomtype.h    d_ticcmd.h    d_mode.h    doomdef.h    m_argv.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    i_sound.h    sounds.h    s_sound.h    d_loop.h    doomstat.h    i_system.h    m_random.h    m_misc.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   stdlib.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   deh_misc.h    doomfeatures.h    limits.h   syslimits.h   limits.h   strings.h   inttypes.h   stdint.h   d_event.h    string.h   posix_string.h   i_timer.h    r_local.h    r_data.h    v_patch.h    net_defs.h    sha1.h    r_segs.h      	��@     �	&zXOf�
�(:
vrh
<�y��f�XZ%Vv+<t>	:LZ(wr��0v�]�<	]J#X<<�<�tY,f
f*K+��	R.X_
	*R[�XY%Wu+<t=	sK[	N�Z�Z	�.� X��igXvLh,t�J<fLgueuj����<�M�rtt/. � x�t�gy<Z�	JY
Jh/	�iJY
J�/	�i.Q	�v��$Yf�=Zd>1fN�0<XKs0.<g�q���ut�-ff<�fs/u�s=Y�=X�H�JR�	JZ=	� JmA JJ		�r�=�=�	\	J* X JOqWJ[	����$Yf�=Z��fJ�f
r>��s=Y�= �J��0	f�%�x�	W�
�(
vHh
	*\Ry�_�	�-�i �ZY	j.f�  ����	'f	XX�	-�t�	<����f�gwf�hf�i	���	���	�	�Lt.�2�vdJ
fh�"<�.]g*g31�vY	F.:X� #Jv<Y	|xX0.1�	f]3�.A[/*.��\r!<u=;=;Y
�Y>�?�
XM�t.�wfu.o. 	iqfJ!k	9iz.u7g0,0,g?GghYgrf�&	<u.vt/?�dlyfm//wfg&'ge==:=(%usKL 	K <Y	< I � - .5�hM7K��ZYX ....� Kw
f	hd!kz<u+?	)hgLh*g�u�&.</?�cfgh��gd1r/&di':e=%/r=(YIg	K<Y	�
KH<-.4�ur1d=d=K=-K>	Y<Y	�I<-..	iX�y5�
X	Kvff�
K
K:iL<m�=�[`J#�<JM
�g<.�J��f�	/	e���=Y	zX�Jztu�X�X..�O7A:!J>[ge=>[]<XK!w.@@ *@� 	iX���u�	\fh�	1Pr� .��h:$X.X'.gtX'.f�z�<L
�#L
�2#ittf��>v:0/hK.0ui�;=Y>t��gY-g.�  w� J�f	.wf	�u<).�%�X[�X[J<�{	=?<�m	=A��Z&#f
��J�Ar�	��/	Zf����gZrhZg
h9=
:>
��X��z
:Z1<.uf<=9v1&tRc�&z�=!�Q!y�<&H0r//&w�	�eN.  =uy.1C<t:u&<KLg&bK�zf=K!N<!8.N&b�X 	A     1	<y�>8v9>,.;#/.s#t=<#-<1X 	`A     ?u
./tf
.=rtJ@pK2o=/@zfK=KI=;K= Y < Y � = X , .1  ..� <�ix| <Y J gE � = XJ , .3 t    r  �      /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed /home/user/.local/share/lemon/sysroot/usr/include/abi-bits  p_maputl.c    stddef.h   m_fixed.h    stdio.h   types.h   stdint.h   m_bbox.h    doomtype.h    d_mode.h    doomdef.h    doomdata.h    d_ticcmd.h    d_loop.h    d_items.h    tables.h    d_think.h    info.h    p_pspr.h    p_mobj.h    r_defs.h    d_player.h    doomstat.h    i_video.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    stdlib.h   alloca.h   feature.h   null.h   size_t.h   wchar_t.h   locale_t.h   posix_stdlib.h   limits.h   syslimits.h   limits.h   seek-whence.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   i_timer.h    net_defs.h    sha1.h    r_local.h    r_data.h    v_patch.h    r_segs.h      	5A     �v4@!.tf	LfLJ�Z<hf%K.-<KA1<jf#K+.J<
.$9uf<w.	J<Y��y�t/t/<K.=./ �LUYJJLYL.nt.>h< j. <<1ue=Z ?+<?  N
�-z>H/;=,�X1	�	X3>H=;/,�X[	�	X3�Ye/2�Ye/�L=.<tLcK\JZYL.w8K?g..g. 1g 0nXX<<<.��=�f?.< </g:/=g z�<<)�t).�.2<f�<s=�#] #.	Y 'J ]J#XJ J� y�!�v*<�YW/*J�2=�/[N��N	�,z#w9/#ru#IK��X�~�Yt (n.?.
�Y�=
Z[/>
�Y
YKLZM#w9/#ru#IK��X�~��...�} w�#K
L"A.t.fLg�gifg f\J�LJYh*Jw\J�LJY[�	< H < f Z g ��<'.t'.N w 
	<fYdL[>�JLYLO[�<H<	f[g��=)�.)t.K<K	YL]"��  �fK�s<Jo  r00�( t J	yf	tJvf:TJ5>.N. 	l X �fK�t<Jt.'tJ J	T|XHJ4. 	t X� v|x<^$MtW YZ	.t2 , J	.	JX<Mo�X<..� j.j<.j<�he.XetX9g�uh�<�h=5=w.=+g8g	
z<	5y<	/]E=z<u<h	IK	LL(
<g-=
��
�J00
;K
t�
�J2
�g�%t%<X[v(
<Y:
g/
 00
W=
L�2
=YZ%J%XXA�z�	l	NfZIYJ0
fh= d< .!.YIY <..-Yt .... �   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_mobj.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_ticcmd.h    z_zone.h    d_mode.h    doomdef.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    i_sound.h    sounds.h    m_cheat.h    st_stuff.h    hu_stuff.h    s_sound.h    d_loop.h    doomstat.h    m_random.h    i_system.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   d_event.h    string.h   posix_string.h   i_timer.h    r_local.h    r_data.h    v_patch.h    net_defs.h    sha1.h    r_segs.h      	�A     �]S]S�)%YW=.Y
LuK
Efo
z<x=g��/�"X[R"u<?�z�ixbw=iZ#+t-/;=>�
Y�'t
<Z
>!��J ... "d>WL�Zt�>.?a�du�/.�<[�=X 	NA     �{gL��M�gcv=@zJg@YZKsg0Y.5+#c=+�$Hv�X�<hA�k�K=Y � k�! X <L&<.1q>-jdhgt[�f�)t3<)<.>	. .	 = eh' . <K	fB�-h X�?<Lu�)=)�=Zv		ff' Xg>Ww!_ !< _ X
�<K��< <<.Mgv[fh?W{.�}.vf�%Ysg"t�l�:vu
�uv<u
�uvKebf��>:J/0,J=2=K<1�M	���tYIZI�:<  ..F.[���X�f�<��ew�%-J	<Oew�Y�!-JfXY����=X<  ..<� xRxt	<�=M
��
HN�
�
�v�w
1z���
'Z
V=t='�h�v�=  -Y  .'"V>0�z���ffvt�	��/�f ����w�X[?[ �  �ptt�����t=M
�
�u�!tf� :�?
0SJ�iGh
'ZW
s=K't�i���J�#p.J<��v�.ZIM	r;?X?Jg!<Xh)�t)q<�g��u����xtu[�tttttvJ.�Z.,ZX	 Jht���K%	�i.�s!g^ ��gW
L[..,\O�<!6Xf� ;�JA" � t���t�9=O+G=>��X=>r"/ Xt�fgggh) gg�.. ��X.Z
�".<
>Y
s=X�<hBz�l/I� YX.�wX.Y
�".<
KY�X�zX<��<
ZYYJ.-YJ.
< =X^
@v<f<gC;.zfl;.=.;=
XK=Y 	 =	Z�U	�	�
 
3)
�f<tX@t<K�
�u
��	X<X<J>rKK/�=��>Yz
z<&O
S0J&<X<=ZJ ..<v.uX
�=-/Z�>0g
�
�>0	g�?0	Y@
Z�
hX>t<K�s>9u"r>�:>�:>...-X  2   {  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_plats.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_ticcmd.h    z_zone.h    d_mode.h    doomdef.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    i_sound.h    sounds.h    s_sound.h    d_loop.h    doomstat.h    i_system.h    m_random.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   d_event.h    string.h   posix_string.h   i_timer.h    r_local.h    r_data.h    v_patch.h    net_defs.h    sha1.h    r_segs.h      	�*A     �2�YYh>�= z<	f#2�Y<'YJZ"=u-� y<	f#2�.�  y<lX�~tufMJY, * J \� ��tvV>2		;=ZEKKK�u>��)Y:u-;4�tYYs=vv2)Wu-4�tY$us=vxu.u�@up0:h2u�?:�Z?r�Xh��<� XXZf  J.0< .?�,J�Y�   v<	fX/�}Xi�Xy<;[	�JXJ\ X�>Is=\	�=uV=�Z�&Z &< Z XvZ>JWs=kZ	J�J].]. �   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_pspr.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_mode.h    doomdef.h    d_event.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    d_ticcmd.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    i_sound.h    sounds.h    s_sound.h    d_loop.h    doomstat.h    m_random.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    deh_misc.h    doomfeatures.h    r_local.h    r_data.h    v_patch.h    net_defs.h    sha1.h    r_segs.h      	�.A     �	B,v�| 	28	xF	$�MJ�1/W�:vh<M;�<kJt_Xvr>yJ�	�<.<u
 u<u+h%g �.#q?/��<�1k1SJh�$�X 	/0A     	
<�X
Z�	W ��i ����
����
���
���
��
��
���
�����$H.�3.' 
?XM�/=/WK�=� 	 $:$0H� 	�1A     tA<u�X[g��. �j,=X ,f<K�h�e[�< t<]�g�=;0;df���Y �. g�hg\�X 	3A     	X 	3A     �xh
w%iJ\�Y
 �r<y /8x/,L� 	�3A      =<XYB<�BJ� 	�3A     �X�HZ/	L�KtY�%.<=ui��LqAf
<�X=JKt[�%.<?o^I/z<B��. .i.[�"3sJJ.<.� ��4 ��@�<.<9!<9XJfY�X9!<9XJfZ�X!W9YtfZ$1�V<�/<:\�.Xj=��h0g��g0	g�i<
 �XYW<JK�X.XX".<0gIYY -X 	�6A      =<XZ�9<9�J�$:$ZH���X#	XtX[<Y�9<9�J�$:$ZH��  � .0.  z4zX.qf.mf�<Y�9<9�J�$:$ZH��   �  < K  t X 2" T < = $ < U$ [ z.# P 9 c/ B G 9 1 � <
.. f.
 KWY<Z6tf��9<9�J�$:$Z����^��.Y. (�#�#�(y	�@�xZt[+:	�7+�:�   X < W <1)t  lf�<
X<X
X�9�gX 	:A     zz	 J�]	tZ�/ t� <�#�. �     �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_saveg.c    stdio.h   stddef.h   dstrings.h    types.h   stdint.h   doomtype.h    deh_main.h    d_ticcmd.h    z_zone.h    m_fixed.h    tables.h    d_mode.h    doomdef.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    p_saveg.h    d_loop.h    doomstat.h    g_game.h    i_system.h    m_misc.h    string.h   stdlib.h   <built-in>    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   d_englsh.h    strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   doomfeatures.h    deh_str.h    sha1.h    d_event.h    r_local.h    posix_string.h   i_timer.h    r_data.h    v_patch.h    net_defs.h    r_segs.h      	t:A     � 	K�	YXX	Z��X /JY=. /JY� /;<� /�X��  �<.X� ��� X�� J� . 	;A     � >[��[������=�yX	 w.3�J> 	 L ,	 0 X0. � 	M�	Z���#X=Z<<1	.MXK�W==W</?=1J	 w.3�J> 	 L V .2. �  ��   �<X� X� X� f^� X� f �~ 	�%Jw��y	�t-�J	uXwY$��	 x*J. @ f	 Y X /	 Y -	 / X0�K�	  f W[v,Y��	  � Wi����'x	 	� W . t	 �  � ;[u�	�-MZ,���   � ;j	�	Z	:=	Y>V".<��#ZX='�"�y.���3�	Z�z�{�f�{.X���~��������������	�V	��Vl�	�Vli+[�	�V	��V	��Vl'�Yf[�������z�����z�����	�}t	Z"	x���<�� ��	����	Z�y�|� �|.X��Xi�XiXiXwXiXiXf� XiXiXiXiXiXiXi	Xt:	�Xt:lX�	Xt:l[+iXi	Xt:	�Xt:	�Xt:l'�YfiXiXiXiXiXiXi�{ X��XiXi�{ X��XiXiXi	�~Zz.	L.J�JXiXiXf�<��X�z�f��� t���x`x.6 t �! / ,5 .! L < Y#  J Y � � � � �3t <�L:Y��	fi	Jv&XY"JY��� uJ* a/ < J.<.Dx`x.6 t � / V5 .$ L g & X g  X K  X K  X K  X K  Y � K   �2t <�
Z:KXK
XK	fh	Ju)XY%XgXKXKXJ wJ* a/ < JX<.<�w ��2 t���Y�v�����~���~������}���}���}������������}���X[�����}����	zz.	Z#-�	@\��}�������}�7 �
 JX/ 	Xy'u�L�X0qXX[Y�Y�u�
<=�u[X?X?X?�~ X�f�~ X�fX?X?X?�~ X�f�~ X�f�~ X�fX?X?X?X?X?X?X?X?Xi�~ X��XiX1XiXiXiXi�~ X��XiXi
Z	L#..t	�	��Xi�~XwXwXwXwXt��~ X�:��Yj8$t/"=�==Y[k<tX]!.% t�J[� ;����Y�z���[���.���Y�z����[��������Y�{��[�����������V���Y�|��[����X���Y�|��[��<X7 � J� XZ�XuY� �!Z�zY�x�<=�x[X?Y.JtMX?X?X?X?X?X?	�X�yX<�#�	/"���[Y�y�<=�y[X?Y.JtMX?X?X?X?X<� �"�\Y�y�<=�y[X?X?Y.JtMX?X?XMX?X<�!�#�\Y�z�<=�z[Y.JtMX?X?X?X?X?X?X?X?X?	�X�zX<� �	/���[Y�z�<=�z[Y.JtMX?X?X?X?#�X�z�<�\Y�{�<=�{[Y.JtMX?X?X?X?$�X�{�<�2Y�{�<=�{[Y.JtMX?X?"�X�{�<��[�� <tX^    �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_setup.c    stdio.h   stddef.h   types.h   stdint.h   z_zone.h    doomtype.h    deh_main.h    m_argv.h    m_fixed.h    m_bbox.h    d_mode.h    doomdef.h    d_ticcmd.h    g_game.h    w_file.h    w_wad.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    i_sound.h    sounds.h    s_sound.h    d_loop.h    doomstat.h    r_data.h    i_system.h    math.h   seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   doomfeatures.h    deh_str.h    sha1.h    i_swap.h    string.h   posix_string.h   i_timer.h    d_event.h    r_local.h    v_patch.h    net_defs.h    r_segs.h      	.QA     � x 6[q'.Mqi[qwZxf . L
  J g
  X t <2/X 	�QA     	�z�	&Y�/u=$T�-lv.o<
t#XuW#.=WgYuV
<u�wq> �t	`gwtuf	Qy<L fg"fg�u$dKJ<K.J	Lh*$<� J�"X20J Xk ]�# <) J J'X/  .-X 	8SA     z 4Ys)<Jg�su[�z.>.g,v f L # V 0 g  f �1/X 	�SA     	z.s<�&XuW&.=Ig�uV<u��u J �  L  8& <* L g . J g  Y � K  X K  J K  J K  K
 � K 1=  .-X 	�TA     x 6$XuW$.=WgYsuZvt .Z
<Y
JgJgJgJK0)XtIeJK0)XtI wf$ .* J J./X 	jUA     x6xX.t<�Y-=%XX..h Z� t  B _X% < J Y  J Y  K W Y   J Z X1uX ..(xfq<�$XuW$.=WgYuV<u��q> �JKJK
JKtXKW=KeK	=	�>K�
K�
	XK�w<<L=\=?JJL=\=?^z.KXLg-2+g, K.% <+ J J:X=  ..IX 	�WA     z.s<z$XuW$.=WgYuV<u�vu J �  L 8+ </ L � ' J �  Y I g  Y � g  X g  X J t X1/  .-X 	�XA      3Y�WuYtmX�<�J�YW<g-8j=u;<uu 
 t.s.�uh r L  # V) . M J � J2�J,u tZLH>�O= x<$ . J J��X�pf f	 N!  ;	 K  . 
J o	 O 3 �	L	�JZ!.J!J.<K	[$J�!.J!J.<KX<5 .�>:Z  h  L : L, < J �,  J �2+J5J&f5<J=)J$J5JJ? �us=- X K  , > # W g   < = >  g e" . f =+  J =  , > ! W g   <  b<* . J <[X � X=3S.=3E=�+����   � � �"��"Z�[�W[x>9YKYK[��0�
<vJY������Y�lz�B*z<<B	Z�	�:�9	Ye	uZ%@	� f�tt.
�%v�

�	@--,	2;;#=0J#<.	K
�	Z�.�		�9[G	[X.� �;�[�	�u-�X 8
f��^�\f.D!YYY 5   !  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_sight.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    doomdef.h    d_ticcmd.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    i_system.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    d_mode.h    d_event.h    r_local.h    r_data.h    v_patch.h    net_defs.h    sha1.h    r_segs.h      	9^A     3<LWM</JtLv
X[Y.L.w9/'?;=
;=	+>Md� �<<)�t).�.2<f�<s=�1	O G[J J(nfKty	JwYX	Jv �Mfa!J<6L=WK�=�[e;	;M�	UYYY�=[	�vyxIK<�&�[	�0<h=	�i��	�ijYXt
<hY.Zfw.<?�	Jw�Y1'
<�N<Q.)<<bXhYLf<	S].  !Ju!d<v;!Jl!zt
K//;@<J
X<=7h3.:h&F/;g/0#q47#eg	>e?*gi	zfg@8ghXi    5  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_spec.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_mode.h    doomdef.h    doomdata.h    d_ticcmd.h    d_loop.h    d_items.h    m_fixed.h    tables.h    d_think.h    info.h    p_pspr.h    p_mobj.h    r_defs.h    d_player.h    doomstat.h    deh_main.h    z_zone.h    m_argv.h    w_file.h    w_wad.h    i_video.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    g_game.h    i_sound.h    sounds.h    s_sound.h    i_system.h    m_misc.h    m_random.h    r_data.h    <built-in>    stdlib.h   alloca.h   feature.h   null.h   size_t.h   wchar_t.h   locale_t.h   posix_stdlib.h   seek-whence.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    net_defs.h    sha1.h    doomfeatures.h    deh_str.h    d_event.h    r_local.h    v_patch.h    r_segs.h      	\bA     ���  .	�KL
9M
	X�t�;Ktx
	XMt�;KtXM
tK';f.>K#
t
=I=
��1<A<+<J1tAJ�Ju 0<@<*<J0t@JH�� "<<J"t)J1Ju 	-iJYM	 0zJB .Z
K�[.X<1	<zJB, ZZ
K�[.X<1<w4z<	�w<	Jw. 	J	hK�	>	[.[\[�.@f.J<3O	M. <	L�5tXJ'zJB, ZZ
K�[<X<1CzJB, 0Z
K�[<X<1<.g� -K<tJ�= yJ	B/ .Z
K�[JX<1<'q
tw[�	�=�X4X�].4X^X^.^.X^.4X4X4�].^.X^X_X^X�]X^XXX��X^��} ]..4�]X^�]X4X4�3X^X^X�3X^X4.X�3��~ ]��4X�3X�g]X3X�<�~ ]�<�~ ]X3X�<�~ ]X3X3.� <� ]X3X].]X]X3..3.X3� <� ].3X3X3X3X4.X4X
.X3X]X]X].X<m ]Y<s ]X3X?[  $~x0�$X<Y3�Yy�Y[[ 
  ?<w�JjgW	<�	�YX.&.Z _i	�
�X	tgg2v�tvg	w \y]  xtR0g/ \ | r z�Z J- J( < JL(5�9.
<=	YhJ</ x. J.,{t y.L�x,X�<.�i<<�Y	0(;�"t.(8<(<8X�1(8�"�� hJ�� Xs	.t<fuJfX��twwJ	�`Xz.of]	JtL	 T���~	�p�	�	�	�	ZJt.X<J�YZ!f�y!�ut.� $=!N=�K#ut�	vX�KuY�M��K#��uKuK�� ��tzBf J	�	�)f��u .�J�\�2O�2�g2�1g2�2y��1�  E* . J� X� .�Jt���)�t'<��<. 5  � ; �  � ;� . �� �   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_switch.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_ticcmd.h    deh_main.h    d_mode.h    doomdef.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    g_game.h    i_sound.h    sounds.h    s_sound.h    d_loop.h    doomstat.h    r_data.h    i_system.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   d_event.h    doomfeatures.h    deh_str.h    sha1.h    string.h   posix_string.h   i_timer.h    r_local.h    v_patch.h    net_defs.h    r_segs.h      	joA     � y ��M�X 0  JZ/<�.g.<n<X<JX=J;u<X�f4�� G�fJ��uggg�K w<fX.X y�Kh!`x.�xXKYzJZd><. <�tLtY7.7X5<)<Z	�4	ZtY4.4X2<&<ZY4<�tY;.;X9<-<Z
Yy C y._  . Lx.	��v
.�J
�U.+tt�
X��y�4�Y\X4X�zz.z.z�4PPz�^z�Y\zzPzzz�^.��
��^����4z�zXzPzX4Xzz.zzz���.���
X�^z��Y g �   G  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_telept.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_mode.h    doomdef.h    doomdata.h    d_ticcmd.h    d_loop.h    d_items.h    m_fixed.h    tables.h    d_think.h    info.h    p_pspr.h    p_mobj.h    r_defs.h    d_player.h    doomstat.h    i_sound.h    sounds.h    s_sound.h    i_video.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    net_defs.h    sha1.h    r_local.h    r_data.h    v_patch.h    r_segs.h      	�tA     -�2Kr.jp0t�:	F� .� � <���
L��KKL�X	`J(t�htY&f?	/�=	t;=	J5�	�����=+�s=
MtJSt� :?�. !   +  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_tick.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    m_fixed.h    tables.h    d_mode.h    doomdef.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    d_ticcmd.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    d_loop.h    doomstat.h    z_zone.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   r_local.h    strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   string.h   posix_string.h   i_timer.h    r_data.h    v_patch.h    net_defs.h    sha1.h    r_segs.h      	vA     .(��
 tK;�u
 �	 (#u�Ji1J>!:=!Kx	YZJ0 	 �wt	 /����. :jYY[g y   ,  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  p_user.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_mode.h    doomdef.h    d_event.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    d_ticcmd.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    d_loop.h    doomstat.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    r_local.h    r_data.h    v_patch.h    net_defs.h    sha1.h    r_segs.h      	wA     7>q�+1#.<XK�=XJ=  .
 vff��V0>�* �� Af=[��h<Z��.x�
Xu	Kw<L#<8f#0:>fK&�.6%7AN)8<@8@�J��J J�<>u<�ZZ   @[<u��v;u;�gZt7 X <Z
<.<0f�>1f
�fK�gu (�yL,vjhiX �K�Z�<&J<u�gL<]*Z:0,1�< T�[g���.�\=�lZ�����<KZ<K$Z<K.Y<�<KZ<KZfK�fK�<LuK
�<H�uM�  l	   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  r_bsp.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_mode.h    doomdef.h    m_fixed.h    m_bbox.h    d_ticcmd.h    d_items.h    tables.h    d_think.h    info.h    p_pspr.h    doomdata.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    r_state.h    r_main.h    r_plane.h    r_things.h    d_loop.h    doomstat.h    i_system.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    d_event.h    net_defs.h    sha1.h    r_data.h    v_patch.h      	�{A     =
�$ y5y<zYYJ0.L.\XYu�?Z	K	IK.��/K2.Z2<#j�[YL<\=3�OXQ��uJ zBz<%S&YJ0.L.R\$1�MYLy/ Y. (�d�g�(x/f9wXu/J�fjibg/;=L1	�0</rJ.J1�	3gg==uwMJw\1tux	�H[tJ{3)\/-Y< �
Z�g-
L�=�%V.%*.VJ%* sWt* =%qz9M<Y;g-/&Xv	u�f1f><L.@-	[0/kJ<Jy.
.[	5ggj.=	=u	wL>YYJ0�J.	� � X. zlfKty	Jsg=KZ*u
Jv�����������.Z=IY0.  hY.Zfv.<?�	Jw�#.$[<9[	�XKiXhYLf. ..  �   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  r_data.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    deh_main.h    d_ticcmd.h    z_zone.h    d_mode.h    w_file.h    w_wad.h    doomdef.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    v_patch.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    d_loop.h    doomstat.h    r_sky.h    i_system.h    m_misc.h    strings.h   <built-in>    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   doomfeatures.h    deh_str.h    sha1.h    i_swap.h    d_event.h    string.h   posix_string.h   i_timer.h    r_local.h    r_data.h    net_defs.h    r_segs.h      	��A     ��JhY0<0/1Y<0K	r<JJ<0.XX0 s.qX�s<J�	���tK� / W��gfJL 1[	�>eW�dK=;W>X�<.<
XI�Y ...-X 	�A     	tX\c<�o�X��"|"xJu���W<Yu  I\�gXfL��<t L L  � / 2 Y I Y2  � < . < . @ �ZJL�2M&su0&V<h80J	.L�#-t#JX<2YX<... $= $v	r="t ="I
�KKX..XZtuZ"�<3 ]$.\�)tW.#XY[r;=J�Z 	 Z Y  � � <0��V=.KX	wUKXZ	XL�V=/X�
4�
-2 L�hYsu!su!su!su!su!su%SvYW=2Ye=	X9JAt<	`Yw<J2X6<<	DY	 J Y% W = X	/Y<	;Y  Y& W = X 6. . M� 3f = $ X t h  J<�Y�wH>WJN	�u�r�+LW	
<vJZW�t.;XuJA����  XL LV=XK! X<=	L.X& y�0 .9 J J.*Xt.t<)YXs=twU>
Y<�.6��	Y r� . f K! - / X10,v  f K  < <0�~XZ,Zr<v�	�.	D	Z1�$t<	L<ZJ	3�f	�<<.�f.|#�9W�\6T.g%f?%qiv,v  �  < </
.$T t.$Y?W�[<q<h%7f.g�su!su v  �0Y �
  !&  t& < g , J u, I g.  � <0. (%��u.!Y�Y�Y�
.	�X0.0K�YYv�f 	-SRx6Z �t<LZ�K	ZJ1=.  
 	iX0.0�J  �n.nX��s=.Z . �  �# � K % � J1� . �0hgW"<��X<2<[!s=.Z . � J �& f K & � K ) � J	.w +L� �f<1
v
:L  X Z  Z � =%  J t � X2�!s=.Z t��",<7 G J4� .�f<. � �Z	� $  f g  �! < � � T f <	.=  �X Y   ~  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  r_draw.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_mode.h    doomdef.h    deh_main.h    d_ticcmd.h    z_zone.h    w_file.h    w_wad.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    v_patch.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    v_video.h    d_loop.h    doomstat.h    i_system.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    doomfeatures.h    deh_str.h    sha1.h    d_event.h    r_local.h    r_data.h    net_defs.h    r_segs.h      	��A     � �w	 Jje	-hI=��&txb"A&a+�
7�
 k %  . y ,% + >0 r < J � h  Y� .�u Jje	-hI=��hwo>"�&b+@)G
1'c&;'�
�=>
 0 . ( . y ,. 99 <( < X �	 J K    vY!.yt'/�����Jjf	-gJ<��&tt&n.
��)t)t�Jt1�l+ciY3w	<������Jkf*jJ<8?��&<)u.'m.&;�'�
�=?)t)t�Jt/+t+t�J	t1�m*ubiYJ�y'Jje	-hI=��&twc"@&b+�
8�
 i 3 . . x -3 + =3 s. <$ J � � g  Y1xD�Jjk�?Y��&t)=1'c&;�'="�a+�
<a=?
 1 3 . . z -3 )$ <3 t. <$ X X � K/ % � �	 � =    uYJ#w]#&"X�'�;K'�t�� t<�&.x(!Wh���gh%ho=@"p;?90g;<
<1%
�� �	     z / A @ v. = Q x. h! @ t X
 �	 > Y �  x(!Wh���ggia=
<"vt;>?)0eCz�<
;1f1�%
� �	     z / A z� = 
J , w. h! @ t X
 J K!  �
 � > Y  [+'..i  K  � <1-�(1t. � . � K  � <� n�	��Y�	Zx�V�Y
v
��t < = I �  ^  x��@*Z"  �% ; = X/�,�  �% e = X/�,�  �  ; = X/�,�  �  e = X1��������.Y
Jt	Z	t.7<J	<<0	 f�%wX%	 j	*�X1
q?
G?�g;<	f=[w	c=
>  � �   q <5X�X    �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  r_main.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    doomdef.h    d_ticcmd.h    d_loop.h    m_fixed.h    m_bbox.h    m_menu.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    r_sky.h    r_data.h    <built-in>    stdlib.h   alloca.h   feature.h   null.h   size_t.h   wchar_t.h   locale_t.h   posix_stdlib.h   math.h   seek-whence.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    d_mode.h    net_defs.h    sha1.h    d_event.h    r_local.h    v_patch.h    r_segs.h      	2�A     � Y=Y=Y=K/ tLcK\JZYL.w8K?g..g. 1g 0nXX<<.�e=ZfC.<(?HI/	/	h.0.9Km�fL[X1/;/+1..Ln.X./;�I=ZfCX e>	?+e/>�y5M\	[XX��<�0	MJX
.�t.�Z[	[�<y�.�0	M�.�t<Xy.	 g,h.X 	w�A     
f/wf	 -.��	J�	0JX.21?1z %.-�?� fX.f. �k74fr<u	Xg	�KZ�L
� 	�J +.t�.t< n< w��K
��1
u#�XZ	Zf w  � pJ�� . �? � ) < � < .4�fY�'
�Kf xJ�g ;g w�pX [�;=<X�&�Xt�t<� ��t �gg'x
<d�Z��/fW�!<� �ei ,> ;g:v<gLH>r<gJuvL
�����
�����Z[&fX&X<g)�bi . K  � < .3 V � L 
  # 0 d
 . . < g   t# /1 J < � t < . 1 f L )  t u) W	 < � X t <1
.#n*�#.?xt1�G1&f?<J�*X#X�v<f ��J!Y��}���~���e�g�� Y�Y�YY��
.	fK	tm �h	=WJu	�
.X1 = -/-Ju(;u��#�eg!8h����hfL�>!,.rx   � ;��gg(![YYY[[�Z[Z[ Q	   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  r_plane.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_ticcmd.h    z_zone.h    d_mode.h    w_file.h    w_wad.h    doomdef.h    doomdata.h    d_loop.h    d_items.h    m_fixed.h    tables.h    d_think.h    info.h    p_pspr.h    p_mobj.h    r_defs.h    d_player.h    doomstat.h    i_video.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    r_sky.h    i_system.h    r_data.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   stdlib.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   d_event.h    string.h   posix_string.h   i_timer.h    net_defs.h    sha1.h    r_local.h    v_patch.h    r_segs.h      	|�A     �  y_���f.Xx$<f�!��!Y!�.�Y��gX���g�Ui��/sK�Jt�g-g<X	>rv\>�
�ugowf...-f 	�A     	hyf% . L  �  � <1t^vf�[zf�iq?��gY� 4z.	�wX&�  tZYg4 T t.��z�?�SK@x.�X .. t�fJX K<w
.|xX=<K"@LzJLx8u+K0l.KM	<J19�J:� Y2J,��Y.<1��X>��<0Xt.	 wt	Jwt	J������� n� ��J�J��l��Y	�g	hLhee,t=Xuf v<	��W=tv��;gxX<fRf0t�JJv  Z $ X	41 Ct t?X  &   q  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  r_segs.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_ticcmd.h    d_mode.h    doomdef.h    doomdata.h    d_loop.h    d_items.h    m_fixed.h    tables.h    d_think.h    info.h    p_pspr.h    p_mobj.h    r_defs.h    d_player.h    doomstat.h    i_video.h    v_patch.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    r_sky.h    i_system.h    r_data.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   stdlib.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   d_event.h    string.h   posix_string.h   i_timer.h    net_defs.h    sha1.h    r_local.h    r_segs.h      	��A     � v
�?(tHIuO18Vuu>)"L)HZHhg
./u
0K
���L:v"+X<;gg�Jh! =/t!;sh \# ���	tYwf pJ t�t	��	03S>t�w#!f#tY2!)=.�!oui.t�
MYt � ' gf f�. Xv� t�< 
  t��?K	>
;K	K
>	ZtY��Y	L�
Y/	K=	LtYyl<� �fs =�kxX=,L>t�,u�J
ffMg9gugXug���]
	�Mf=�KYLZg9gugXug(�.�
	�M
��8=�K>Zg9gugXvg�<�	�t�#�~f�fg
��x�tJ�XXwt�Mcw%�g%f]1�;/!�2.!u<=,K�rci	{yf=Ko=�	WtfMZA<'h:�rK �!IfXO+t	�oI=[-��,�+-,=+-,u	ipg��[)!J���h��15�Mh�w�+)9��vLuZ
L�-JZKh
LKxLH�uZH�u(%=?%c(;@pu%Xw/XZxbL(xbZ
(K[��[-%X�u	����M0(X�hyJgi�>��>�K0euJ�+�;ffhh�Lu.0!�!I<=�dh��/&t�g%�%z�l0v#<*H	>*:Xh	Y./g0	K���"tfM�YJ��ids�Y"t�/Ig"Z ��Y%t�/Ig%#X>#�vhgs?cg0#t�K!��X�f�"t�K ��X���v��v\t(f�v5"fX5�+..Y!u��t+f�v3 f<3�)..Y$u��  � <Z=s= <Z=s=	�X� �   �  �      /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  r_sky.c    m_fixed.h    stddef.h   stdio.h   types.h   stdint.h   doomtype.h    doomdef.h    d_think.h    tables.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    d_items.h    p_pspr.h    d_ticcmd.h    r_state.h    r_sky.h    r_data.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    d_mode.h    v_patch.h    net_defs.h    sha1.h      	+�A     /� �   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  r_things.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    deh_main.h    d_mode.h    doomdef.h    d_ticcmd.h    z_zone.h    w_file.h    w_wad.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    v_patch.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    d_loop.h    doomstat.h    r_segs.h    i_system.h    strings.h   seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   stdlib.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   doomfeatures.h    deh_str.h    sha1.h    string.h   posix_string.h   i_timer.h    i_swap.h    d_event.h    r_local.h    r_data.h    net_defs.h      	6�A     � i�<Xw�h�[K?J�[$Mt+�   �  � 9	�K?NF�t��#*J#uI*<�%�<JX=gJ0<Jho�.lt�l. Dd.JZrve=OJ X�Y�z<BT�uL �t�<	�LY	�=>��X���JZ"I>�= nX <��JZ�[
0<
:h  fZ�pJ<tfh. Dg
���+ nt <�	v	r<K��Lt�<[X �   3  � :�X 	�A     
�	 t��	\ kh<�&-g&I/;<ggLt q=;g:hJK��K ��8%<!-%K!-u%kh1	JX[g.  y5yX�f�Jv[
�<v
*v
�u+�x"fg;? =p/
gH1"c�" X> :v f�t, . JY �   <	 W >- wX6 f J.�. .
<b
?
cg
L
,vY�=Z?��yJZ�0Y�/Y1	tJ�J��LH>,JvXg�4%�JLw�JX=gf3gfNt=-Kt�M�u-gX1�?.jZjzt=t=uuuJ=J= g;=�=-f J < =  � vu$-f=2u?<Y) <J=M�
�t
]q	t"�S0f�L�
 f\t >!�f/
��� J Y1 � J0  'sX�Xw!J0!:>,JvXK�1	J9wf%�JL#YMF=htKt�M�uegX8�?.jB�V�B9Ju9;KKeK- J = � K  . L fZg$tfjK�Y) XXL
Tt,J<uM
�t
]Ji��[��...(z't<$J1<�f/
���x���/yW�
yZ  #vV�yX> [ Z  K s K  J1u Oy.�K \/�� Z	Y	Z <Z	J�- : J 6  < tJ . =  u  s �  =  u s K 0
 w.	� t K  � � <3tJ ��<�J�g�19=v<�XO	�K�XJ>�>�>.�X ?��%��<0
< [Y�"��<0
< [Z�%���"��<) �. J� X �L����<1�;� ..-X 	��A     
$Z��v. t�
J	.u) � J��Y  �	   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  sha1.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    sha1.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   stdlib.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   string.h   posix_string.h   assert.h   i_swap.h    strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h     	��A     7%)]K<K<K<K<	P Z / d L =  g  g 	 a X�Y��G>>Yo�KN��u.X�����<�<�����rt�������� ����������=>:0�9X�Vt�/<;�X=W��;f<�*<g;��f<f� .�<=-�֬fX�<�t.�XX�K;t�f�X.�.t��<t�<�.t �� fX�� fX���V��>:�Vf�:<��<V�<��=W�fuZ�;�Vh:fJ�h.�J�,�J=etf�gW�=/-I�K=H=-Z;;�=-�Iusv��=-<Y1Tus=|wX���=;M�-�:L:X�.J�W�ff�<fJJ<g�K;=;�ffYW�Wg;g;K;=<W��fJ�. �.�t�X�<ɝ/?Tt%-<t�t<X>V�:�W�/.�X�<.�J<J<X<��.J�.��X�X��<.J.t��f�It�uWg;K;��.J<XX�<�XXX��.t.J�t�JJJ.�JX.J��Y�t�V�<.J!YV���;g�JY;xF�uWtJX�I��Xg-/I?9g>G�Z,Z,���t.<�KIJtKW�<=;��X�Ȑ��<��f�fJ��f�fJ��f.=;.KT<�<YCxX/4yJ=]zJ<@T<�?U<@I>:==KJ�~��zt>��� �;=[JY>9u.� L X J Y # <' ; = < <g�<q.�fh?GYu=.zJ ` X J Y  f t J/ ��*$<*t>	G-=>/>	�	;=	0?<U\JYfzJYfu(��HhAz<LFN�J=X=X=X=?c?�. .?znSO�[(=tJ(<fX  S   M  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  i_sound.h    sounds.h    sounds.c    stdlib.h   alloca.h   feature.h   null.h   stddef.h   size_t.h   wchar_t.h   locale_t.h   posix_stdlib.h   doomtype.h    strings.h   inttypes.h   stdint.h   stdint.h   types.h   limits.h   syslimits.h   limits.h       �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  statdump.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    doomdef.h    d_items.h    m_fixed.h    tables.h    d_think.h    info.h    d_player.h    m_argv.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   stdlib.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   i_timer.h    d_mode.h    p_pspr.h    p_mobj.h    doomdata.h    d_ticcmd.h    net_defs.h    sha1.h    statdump.h      	]�A     � 	=XX9 J# f	Z	<�,	vd	fZ #/ A   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  st_lib.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    deh_main.h    doomdef.h    z_zone.h    v_patch.h    v_video.h    d_ticcmd.h    w_file.h    w_wad.h    m_cheat.h    st_stuff.h    m_fixed.h    d_think.h    tables.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    st_lib.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    i_system.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   ctype.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   doomfeatures.h    deh_str.h    sha1.h    string.h   posix_string.h   i_timer.h    d_mode.h    i_swap.h    d_event.h    r_local.h    r_data.h    net_defs.h    r_segs.h      	��A     3!�u.
G/
=u=KK
K 
IK
8>
�K
YLZ
gWZ
gWX?2t>�X�X���M<KJ3!s=!< !fJ!J<� JnY�IK.J.-YfJ..(	J XY �	
� �X/
=�KK
J� 
K	 � J JYt.ZY . 	{�A     
/
=uKK
K(	J$ � J$ J. .: �z��xRZJ=;�KU=J/	��XZ�"J"X<�f>Xf 
/
=uKK
K(	J�!Jy�	�w	.K;=IYKV/��JY�u<w�	Ju <>f?. ...< �   ]  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  st_stuff.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_ticcmd.h    d_event.h    i_video.h    z_zone.h    d_mode.h    w_file.h    w_wad.h    deh_main.h    doomdef.h    g_game.h    m_cheat.h    st_stuff.h    m_fixed.h    d_think.h    tables.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    v_patch.h    st_lib.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    am_map.h    i_sound.h    sounds.h    s_sound.h    v_video.h    d_loop.h    doomstat.h    dstrings.h    m_random.h    m_misc.h    p_inter.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   i_system.h    strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   doomfeatures.h    deh_str.h    sha1.h    deh_misc.h    string.h   posix_string.h   i_timer.h    doomkeys.h    r_local.h    r_data.h    net_defs.h    r_segs.h    d_englsh.h      	0�A     �	 =XX= � w 	 � � X	 Y z�f� 	 u � qm� 	 � �  � x�f�x.K��i< >$ V > Y �  l	 u � 	 u � 	 u � 	 u � # l. .	 Y � j���X J< =Yu �z 	�	$���	0Z$m	.Y>Zi�
X h� �����~�
�L!;g0<Y�u���Lu�   � Ijv�L[�Lu�   � Ijy�MZ[��u��_� ��!&<><[	f$<><YhO���d�R":h/v��B�� .<L�g	�g�v  u<f
�Li�L!t�#u��	L*�	G$ "�
�Z<<Iy=A
�
b_
N
Y[
Y[
K�
Y�2ue�Xt.At��$A.Y.eA<<�
tx(f�th���fXZ�2.t�eX Fn	M��&X�9GX�
t�t�<��	�Z�&X-�AXtfM/W/k/��NZ�Z�f�
t�	�Z��&X\��&X��
t�	fY�.��Y�&��lX��t�h���.�8XY��8.%��h1y'& �[
��#<�#hVv/t 7	f[m�irt [q� ��x.g+JKL. 7	�
i1"gXgYt�3yt	 	:hM).)X<.^L<
X>i
.1fL
�>i
<1
>Vu
u	X!�>��g>f�><N[ #x � J w + i  r � , � Z  � ���  ������v X 	��A     "�[Z]xV$" J � g!  � < i [  �  
0
� .�!�g
.�2t����u�ts�v 1  �j_
wt3�%!�ZX.	 <k..jF	�wc?�i	�' L  , �  � , v . : u ; � �
f	(%1%%%444	44444t�$���m<"�ZYY�.!Y"u �     �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  s_sound.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    i_sound.h    d_ticcmd.h    d_mode.h    doomdef.h    doomdata.h    d_loop.h    d_items.h    m_fixed.h    tables.h    d_think.h    info.h    p_pspr.h    p_mobj.h    r_defs.h    d_player.h    doomstat.h    sounds.h    s_sound.h    m_argv.h    i_video.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    p_local.h    p_spec.h    w_file.h    w_wad.h    z_zone.h    i_system.h    m_misc.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   stdlib.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   d_event.h    doomfeatures.h    deh_str.h    string.h   posix_string.h   i_timer.h    net_defs.h    sha1.h    m_random.h    r_local.h    r_data.h    v_patch.h    r_segs.h      	��A     �!Y\$tv	j<XL	�

<	=v � x�#<KI#/;	<�	f�1<1J7J.0�,&.<�J	L.	2M?=Xw�M	0
L	�(�#->(W6.<=:	_%Y%W3.<=:3�t�~ � .	L$ fh.+ T .n� x	tw	��<	Z.Xw�	v	�	�fLQ3 X J	Z	%0
�s�	�	���~<�<[�~�	ZjXh�+w.<ff<]�<3�	:LJ'tJ	�R�<	� t�J	� J�t?=L�<�EA	0�?�tX=�C �	�	#Y�? �	�	#Y�Cx
�v.RZ  �	h	�	LZ�MiV�K0�OL PJ�%:P�6.X<\X<.? /	Z�\/X 	h�A      /	Z�[g �| ?U?U#Zuy1f+w 	 L  t �2�	 30  � ��YY�X\	�#�	[Y��u�	��<x�  Y ��<	Z.qt	.X2<��[	h��?�:L�-K�uX �| z&z. P	��ht<3hr�:	4	fZ+..<.2!.fIYX 	��A     �t  �   �  �      /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  tables.c    types.h   stdint.h   doomtype.h    m_fixed.h    tables.h    strings.h   size_t.h   stddef.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h     	��A     )V	�!t<2T	0� 4     �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  v_video.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    i_video.h    v_patch.h    v_video.h    w_file.h    w_wad.h    z_zone.h    m_misc.h    i_system.h    m_bbox.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   math.h   d_ticcmd.h    strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   d_event.h    deh_str.h    doomfeatures.h    i_swap.h    m_fixed.h    d_mode.h    config.h      	��A     � �	�.z	B.z	BXz	&Y	�  .	,X ��YK�K�K�J	vXx�&.f ;&g ;.=
<'s	<Y 	 Z �	 s /   p <4f.... u(w
	tJ
/I/1q?_�	o.��K�J	v�1c�L*-<<v J	L/X	?<Z.�+=Zt�K0:JX.<1.	<w
	tJ
/I/1q?_	o.��J=�J.	v��c�	Z*-<�v J	Z/J	?<Z.�+=Zt�K0:JX.<i.
<X 	�A     
z
zJ
/I/.Y<=�J.	vXwhY+-<<v J	Z1X	@<L/uHK=.Z%4<Kf,;2<"<2t"<Jg0<JX.<1.	<z
zJ
/I/0r>^hY+-<<v	x..�f< R	Z1X	@<L/uVK=<h* <K=3d&<<&t<Jg0<JX1.	<z
zJ
/I/.Y<=�J.	vXwhY+-<<v J	Z1X	@<L/uHK=.Z%4<Kf,;2<"<2t"<Jg0<JX.<1.	<y
�J
/I/.Y</�J.	vXw-fwY*&=-�8=W=> �	Z1X	@<L/�FK=Z&#X.t#tJK�Yt1<JX.<1.<{!�u	.!�u6<2YK�<vXx0d�*<
<v<h�s.=0  ...#'+f'<+<	<t> . J	 2 L  J <	 1  wt ..#'+f>',+<	<v 	 L  < <0#'+f>',+<	<v 	 L  �	 = 0# =;�Y��Y�	.=�/&%u%�( zzz<4zJBzX^z.^z�J^X	XkX>zXKG�\zJYY/KY
pg1 .ZX�.<1=XJ<<3= 0 
 J J ;�ue=ZI=  ..IX 	6�A     � 	mXm.	J�� F .
X	���:�X &u.u��uXJY�KY�=Ye=Y�=Y�=]. � �. � � �
����f	P0/�	K3<	fw�	Xw�2OZ	,	Z�><�^H�ZZ...,ZX<... i   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  wi_stuff.c    stdio.h   stddef.h   types.h   stdint.h   z_zone.h    doomtype.h    deh_main.h    d_ticcmd.h    d_event.h    d_mode.h    w_file.h    w_wad.h    doomdef.h    g_game.h    m_fixed.h    tables.h    d_think.h    doomdata.h    info.h    p_mobj.h    r_defs.h    d_player.h    i_video.h    v_patch.h    d_items.h    p_pspr.h    r_state.h    r_main.h    r_bsp.h    r_plane.h    r_things.h    r_draw.h    i_sound.h    sounds.h    s_sound.h    d_loop.h    doomstat.h    v_video.h    wi_stuff.h    m_misc.h    m_random.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   doomfeatures.h    deh_str.h    sha1.h    i_swap.h    i_system.h    string.h   posix_string.h   i_timer.h    r_local.h    r_data.h    net_defs.h    r_segs.h      	hB     � =XX= �~ 3 � � u . .-.� XX " . +	m���	t v � t��;=J <�����J<f< X	 u � pn������	�M	 ����k.�������� 	 � � f	 Y x�ff	Z
Z�! X^]�X"� =Yu �u �A�  �	�"t	X"X	.$J"<	J$2t	Zr.2<<$>"<	J
�	5	�Zz$T$T$t .<J%.tX�J.<< ><Jj *t 	B     
ttf"�<uq"XgJ?!�X<>	XA� JnX"Jg<?!�J<>	JA�w�t�ty�
f���	+wK�)Xg
Y(�2X&J�
Y�<<..<#�ty�
t�<��fZ#X�%u2	�Zu#X-X!JQ��<g
 X&=<<<XX#�tyX
<���JK�<.   �
tKLn3X	!-/R	A��.k.XX.Zs=< �.<J�Jtt2Y<t��J'I\tjY�  -X }�xR�\d
=�
>:
K#X�K	 X < <K�fktH>H.X  ..<
 ��	�""Z�[4��	�\!Z
� ��0<�g1A[Z	�ti�tZh<\*< X [  . K s / X1	tg��@�M�\
yX5��J 7fO �+���1�� Hj� xJf^y'Z ���	��	#
�"Jt HjX� x<ftY�f���	��	�
�&<JZGKNYh.�hf p�fZY�.S�� c<!�ZtY
�Z��	�s Zu 
[L���3x&�bX l.([Y[/X/��/� xY[���&b�&< x/��/< x	��#��#t x�,f�,t  t    a<#��	Jy�2� �  Em �  q<ft.C(8�����=�.:���
X� y<
f�h^y'Z ��1{
xu<�
	y�	�%,JX�%,XX�'.XX�	Y��< vJf��fZ��6t�	�"�Hh*1f	XK�X vJ
�Z�
�6t�	�"�Ig*1f	XK�X wJfV�
^�� �8t�	�#�Hh,3f	XK�X vJf�.��
�Z�z�f	�"�:�"	XY�f v<fZXu
�Z��	�s Zu 
[L���3�rX$
t>[Z[t��'J<�t��)t<�t��)t<��t��< &f<xt5yfXL�u;�Y�<v���<v�Y.0�2s�X0X2s�X1X�3q��J m<�<J]���1!������\"Z ��y.)s�"�)JJg")JJg$+JJg�g=W
<gY�fZv��3tt'�.JJ�g
2Zv��3tt'�.JJ�g�
�Zv��5t t)�0JJ�g
3Z��!hV>t!�g!-/
>dh
>
rhfL	dh	
{Z��	�r Zt 
[L���1$T2�<Z[?vJZZYL/"/"YLtZY�[+[<#aOXt��	Jhv�v1�	hv�v1�< m< f�&	0�Mu�1�Z.vX �  r.Y
 �  s Yt \x `�.!���3	Tx^�
�wXu	.�x��..sX�Y
�Z\_$?	gJt�gG	��v/vgvgv�
.YX#!YZ�
Y�Z /   +  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  w_checksum.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    sha1.h    w_file.h    w_wad.h    stdlib.h   m_misc.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   string.h   posix_string.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   w_checksum.h    d_mode.h      	\B     � �u.�\XZ� 	 �1  k.1 �	 J gt   � X �$  `J  v�	Z<	�Gs��v&Z	Xo.Y�Y�XX�	    �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  w_file.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    m_argv.h    w_file.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   config.h    strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h     	^B     5w 
	<XZ		�	w . 	yB     << 	B     <<  u   �  �      /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix  w_main.c    stddef.h   types.h   stdint.h   doomtype.h    m_argv.h    stdio.h   w_file.h    w_wad.h    d_iwad.h    doomfeatures.h    d_mode.h    strings.h   size_t.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   w_main.h    w_merge.h    seek-whence.h   feature.h   null.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   z_zone.h      	�B     ��~	�.�~�	�.u�~�.�.  � �ZZV>XY�xX. �   }  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  w_wad.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_mode.h    i_video.h    z_zone.h    w_file.h    w_wad.h    d_iwad.h    i_system.h    stdlib.h   strings.h   m_misc.h    string.h   ctype.h   seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   posix_string.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   config.h    i_swap.h    d_ticcmd.h    d_event.h      	�B     � y� [ X	 Z.  X X X ,l<<8 sX>Z�Y
[f	<X,h-<	XX	J�x._y<=g(OS]Y	]><M<L�
K
s=	v�	>YN�� �u��Zt,�Z<�	Z!�	JZJZ�	%tXZ0<�/�#ft<�Y� �<�� �Ju� >  Z  I K  �# xJ < M =  K � =  Z  1�t	ZY��`
tzlztz	Z	Z%L<	 XZ�Lt> � J .	.	�L<$H..=f
 	iX0	L�[J ( /�twJ�
.b�0.t[fvZ	0<L�\/ -X��.t[
t{�	\/J<
0J	\l<�J�;K	�MX ..(JKXKIt ?�tw
JvJ	z�	� #!Y� Jyt	Z\f	L2<	w+	Ye<	u�	 t Z +  � �(  X t K  < .�	�'fZ�Lt< xJf�    �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  z_zone.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    i_system.h    <built-in>    z_zone.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   d_ticcmd.h    strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   d_event.h      	�#B     � LGIN!LJJOx.u:v=(N�OzJuF1"s<N!LFKuJMv"=_$Lz^�Xv' f J[xFu�Fv	1	YJ	K	Ltgff<K	i	KJ	K	LtgL    x6Dp
`x<
tNl
<�J�J>	[	�<Z\J_K�KJ3M* f# .\>	[<	=	0G	u	�	K	K	L	K?��KHL	Z@�v. .... pf2 K �]9MUi�J pXX  <q�U#.��JXYMtJJ^<<Y�Jg� f�5m�L.  .'#U[0��tJJ^<<Y�Jg� f�5n�LX. (q#LtJJ^<<Y�Jg�* f Jg5q�L. 	 3	�.<Xw X	u#=. ..#�	�XwKK. (
r0K I	\<�+J5#� �   �  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  w_file_stdc.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    w_file.h    z_zone.h    m_misc.h    seek-whence.h   feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h     	)B     � x6x.|x. DJ\w� +X 	Q)B     f AJY=X 	g)B     c$T2X>._:s=�YI==< s   h  �      /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed  i_input.c    stdio.h   stddef.h   types.h   stdint.h   doomtype.h    d_event.h    i_video.h    i_scale.h    m_argv.h    m_config.h    m_fixed.h    tables.h    v_video.h    w_file.h    w_wad.h    doomgeneric.h    stdlib.h   alloca.h   feature.h   null.h   size_t.h   wchar_t.h   locale_t.h   posix_stdlib.h   ctype.h   math.h   string.h   posix_string.h   fcntl.h   abi.h   fcntl.h   seek-whence.h   mode_t.h   off_t.h   pid_t.h   ssize_t.h   stdarg.h   posix_stdio.h   config.h    deh_str.h    doomfeatures.h    strings.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   doomkeys.h    i_joystick.h    i_system.h    d_ticcmd.h    i_swap.h    i_timer.h    m_misc.h    v_patch.h    d_mode.h    z_zone.h      	�)B     �K	�	�g�	k.PSyU	@f	NP0t��� KHo	0L<t22&LL��� R�L�[ -	     �      /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include-fixed /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix /home/user/.local/share/lemon/sysroot/usr/include/sys /home/user/.local/share/lemon/sysroot/usr/include/bits/ansi  i_video.c    stddef.h   types.h   stdint.h   doomtype.h    v_video.h    m_argv.h    stdio.h   doomdef.h    d_main.h    i_video.h    z_zone.h    m_fixed.h    tables.h    doomgeneric.h    stdlib.h   <built-in>    config.h    strings.h   size_t.h   inttypes.h   stdint.h   limits.h   syslimits.h   limits.h   v_patch.h    d_event.h    seek-whence.h   feature.h   null.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   string.h   posix_string.h   i_timer.h    d_mode.h    doomkeys.h    stdbool.h   alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   fcntl.h   abi.h   fcntl.h   mode_t.h   pid_t.h   types.h   id_t.h   uid_t.h   gid_t.h   dev_t.h   ino_t.h   blksize_t.h   blkcnt_t.h   nlink_t.h   time_t.h   suseconds_t.h   fsblkcnt_t.h   fsfilcnt_t.h     	g*B     � �	Z�	�$=<;=;=>-�	Z<2#"?czf	("Y�	�YW?	�"�?��",�?e	=f	>	 < �0 = � < Y"  � . . K  <& + <	 ^  p<�1o�� ovvS�w��v.��[B�	�	Kt.	�W	gL f	w U/ s	/�	�y-�uO���v\!�u	ffv!
�ku1zt!@.Z�T>Z:LX[[	 < �  	<& v� 
< �I 3 �N � . <	0t.^fv,^td<<0. .J-_� +r+0	 �  s /	 �+  J	 �+  J	 �+  J ��%foJ<.s<Xu<Z,
W
.;8	f	4 pJ .�tX 	�.B     #< A     �      /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include  doomgeneric.c    types.h   stdint.h   doomgeneric.h    <built-in>    stdint.h     	�.B     !�v/ �   �  �      /home/user/.local/share/lemon/sysroot/usr/include/gfx/window /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/lemon /home/user/.local/share/lemon/sysroot/usr/include/gfx /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0 /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/bits /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/x86_64-lemon/bits /home/user/.local/share/lemon/sysroot/usr/include/abi-bits /home/user/.local/share/lemon/sysroot/usr/include/bits/posix  doomgeneric_lemon.cpp    window.h   stdio.h   stddef.h   types.h   stdint.h   types.h   surface.h   graphics.h   cstdlib   std_abs.h   c++config.h 	  stdlib.h   stdlib.h   list.h   ipc.h   doomgeneric.h    string.h   ctype.h   <built-in>    seek-whence.h 
  feature.h   null.h   size_t.h   ssize_t.h   stdarg.h   posix_stdio.h   off_t.h   stdint.h   syscall.h   widgets.h   fb.h   posix_string.h   os_defines.h 	  cpu_defines.h 	  alloca.h   wchar_t.h   locale_t.h   posix_stdlib.h   keyboard.h   doomkeys.h      	/B     � o X/W#$.Yd.X.X1Xn.X4X+X4X!$d*<<3!*:�/�#$�Z�	�vu1K�YY��/�	y#tu�[3-!3f�/1-#g�K1
j*�/-��Y0
X#!t�	JY>Z  	@     ���� �    �   �      ../src /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include ../include/lemon  ipc.cpp   types.h   stdint.h   ipc.h    , 	1B     ��	�K2>������ �   Y  �      ../src/gfx /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include ../include/gfx ../include/lemon /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0 /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/bits /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/x86_64-lemon/bits  graphics.cpp   types.h   stdint.h   surface.h   fb.h   graphics.h   stddef.h   cstdlib   std_abs.h   c++config.h 	  stdlib.h   stdlib.h   <built-in>     ? 	�1B     4� Y�	V2 ?0=tY Y�	V5��� Y�V	x. <0=t+ X tY	g[��t. X tY��#u	��E1,���tgXuXuJ�Xv�K01�!<b<, J9 <G <; <# .R J` <I <k Jx <� <z <b . J t 
Y>��X t f . =E0&�h>(ggwgg)w5�0t;.f�� t% �5 � tK0�$t<A.�5tI J5 t X <	 >g:f/�� w��]>8�J/<J&JJ�U>��
XL%K(�.<�4�6<%=��vu t �, � t� t �- � t.�$� f2t�Z JP �L f_ Xb X9 �� J� �| f� X� Xi ��(�-tJ><C�J<Y2�.f@t��@f<@/6�2fEXHX���H< <@/6�2fEXHX���H< <�F  � g t w<�o>�ggwggw t$ �4 � t� �� X� J� t� J� t� J� �� J� t� � Jn <| Xq J� t� J~ t� Jn �� J� tc � J6 JD X9 JS tH JF tU J6 �` J\ t+ � J .�_>)+w>�ggwggw#�*t6 J* t X < > t% �5 � t� �� X� J� t� J� t� J� �� J� t� � Jn <| Xq J� t� J~ t� Jn �� J� tc � J5 JC X8 JR tG JE tT J5 �` J\ t* � J ,�D>
= t! t. �> t5 <! J �)<"t8.?tG JV t? < f t{ = f[ .k �e tp Jb f  J> �4 t, J6 fP <G <' � < ��V>#%6<%<@.FtN Jd tF < f	 <$ =7 <& <A .H tP Jg tH < f	 < = <2 X9 tA JP t9 < f	 <
 = t, �< t3 < J� Y f[ .w �g < Xy t� <� f� <� f  t> �4 t, J6 fP <G <' � < ��O>�
� t! t. �> t5 <! J� t! t. �= t4 <! J�tf"t$<KuEtQfTt�<"Xt(<5X,<6JT�8.2I  �� )   �  �      ../src/gfx/window ../include/gfx/window ../include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include ../include/lemon ../include/gfx /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0 /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/bits /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/x86_64-lemon/bits  window.cpp   window.h   list.h   types.h   stdint.h   types.h   surface.h   graphics.h   stddef.h   cstdlib 	  std_abs.h 
  c++config.h   stdlib.h   stdlib.h 	  <built-in>     , 	�>B     
7�"	�KZ>R�	�K%><�"/L@��'L�M/0�!�/	��?�=�">�LL	;K v�	�J	 XK��>��$L�!��Y��O+��L>�+��<�
&, t � �.   f -
j�Y���7>
�, t �,�1�fK0'���x.�8>
��K&�;�2��-�"	�Y;0�
��K&�=�4��yX2 t �,�1�fK,#��y.�,>�/  	�DB     �*  	�DB     �t  	vEB     �  	�EB     ����  	�EB     	 � t J /  	�EB     � 
�u  	 FB     � �t J t! X t7 X> th�/ t+ �$ t; X/ tF X �h�  	�FB     � �  	�FB     �  	�FB     )�#���tY��Y����  	�GB     � �t J tZ��/ t+ �$ t; X/ tF X �h�t! X �0 XF t' �K�! X t0 XF �' t=" f tut�tf% J ��
�K �    *   �       ../src/gfx/sse2.asm      	�HB     !>==ALLKK0=!#!>==?LLKK0=!#!>>K0YLKYKYKYMKL1="#!>==>K0YLKYMKL1="    �  �      ../src /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0 /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/bits /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/x86_64-lemon/bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include  runtime.cpp   cstdlib   std_abs.h   c++config.h   stddef.h   stdlib.h   stdlib.h   <built-in>      	�IB     �u��2�u��2��@��@��@��            __MLIBC_INT_FAST32_C(x) __MLIBC_INT64_C(x) PRIiLEAST32 "i" __SIG_ATOMIC_MAX__ 0x7fffffff __FLT64_HAS_QUIET_NAN__ 1 _GCC_NEXT_LIMITS_H INTPTR_MIN __MLIBC_INTPTR_MIN WCHAR_MIN __MLIBC_WCHAR_MIN __LDBL_MAX__ 1.18973149535723176502126385303097021e+4932L __DBL_DECIMAL_DIG__ 17 __FLT64_MAX_EXP__ 1024 __FLT_MIN_10_EXP__ (-37) _IOLBF 2 __FLT64X_EPSILON__ 1.08420217248550443400745280086994171e-19F64x __FLT32X_MAX_EXP__ 1024 __GCC_ATOMIC_TEST_AND_SET_TRUEVAL 1 __DEC64_EPSILON__ 1E-15DD __DBL_DENORM_MIN__ ((double)4.94065645841246544176568792868221372e-324L) __io_mode __INTPTR_MAX__ 0x7fffffffffffffffL __MLIBC_INT64_C(x) __INT64_C(x) __FLT32_MANT_DIG__ 24 LINUX 1 UINT8_MAX __MLIBC_UINT8_MAX __FLT128_MANT_DIG__ 113 INT8_MAX __MLIBC_INT8_MAX stderr FOPEN_MAX 1024 __buffer_size __FLT32X_DECIMAL_DIG__ 17 __k8__ 1 __DBL_MIN_EXP__ (-1021) __INT_FAST64_MAX__ 0x7fffffffffffffffL PRIdLEAST16 "d" __GCC_ATOMIC_CHAR16_T_LOCK_FREE 2 __FLT32X_MAX__ 1.79769313486231570814527423731704357e+308F32x __SIZEOF_WINT_T__ 4 __UINTPTR_MAX__ 0xffffffffffffffffUL PRIuFAST64 "lu" PRIXMAX "lX" INT_LEAST32_MAX __MLIBC_INT32_MAX PRIXFAST8 "X" EOF (-1) __GNUC_MINOR__ 2 _GCC_SIZE_T  __CHAR32_TYPE__ unsigned int i_main.c __need_NULL  __FLT64_MIN__ 2.22507385850720138309023271733240406e-308F64 __LONG_LONG_WIDTH__ 64 __GCC_HAVE_SYNC_COMPARE_AND_SWAP_8 1 __FLT_DENORM_MIN__ 1.40129846432481707092372958328991613e-45F __CHAR16_TYPE__ short unsigned int __MLIBC_INT32_MIN (-__MLIBC_INT32_MAX - 1) __SIZEOF_SIZE_T__ 8 MLIBC_POSIX_STDIO_H  UINT64_C(x) __MLIBC_UINT64_C(x) __ORDER_BIG_ENDIAN__ 4321 __GNUC__ 8 __SIZE_T  FILENAME_MAX 256 __UINT64_C(c) c ## UL __DBL_MANT_DIG__ 53 __FLT_HAS_QUIET_NAN__ 1 __FLT32_MAX__ 3.40282346638528859811704183484516925e+38F32 __MLIBC_UINT_FAST8_MAX __MLIBC_UINT8_MAX __INT_MAX__ 0x7fffffff __ATOMIC_RELEASE 3 SIG_ATOMIC_MIN __MLIBC_SIG_ATOMIC_MIN _IOFBF 1 __MLIBC_INT8_MIN (-__MLIBC_INT8_MAX - 1) __INT16_TYPE__ short int __DEC32_EPSILON__ 1E-6DF __OPTIMIZE__ 1 __LDBL_DIG__ 18 __FLT64X_MAX_EXP__ 16384 __ATOMIC_SEQ_CST 5 PRIiFAST32 "li" __MLIBC_SIG_ATOMIC_MAX __SIG_ATOMIC_MAX__ WINT_MIN __MLIBC_WINT_MIN __SIZEOF_SHORT__ 2 __UINT64_TYPE__ long unsigned int __INT_FAST32_MAX__ 0x7fffffffffffffffL __INT_LEAST8_TYPE__ signed char PRIxLEAST32 "x" __UINT_LEAST32_TYPE__ unsigned int __MLIBC_INT_FAST16_MIN __MLIBC_INT64_MIN __UINT_FAST32_TYPE__ long unsigned int __BYTE_ORDER__ __ORDER_LITTLE_ENDIAN__ __LDBL_MIN__ 3.36210314311209350626267781732175260e-4932L __FLT32_MIN_10_EXP__ (-37) __DBL_HAS_DENORM__ 1 __INT_LEAST64_TYPE__ long int __WCHAR_MIN__ (-__WCHAR_MAX__ - 1) __STDC_UTF_32__ 1 __INT_LEAST16_MAX__ 0x7fff __FLT32_HAS_DENORM__ 1 __SCHAR_MAX__ 0x7f PRIiMAX "li" __MLIBC_INTMAX_MIN (-__INTMAX_MAX__ - 1) __FLT64_DIG__ 15 __ATOMIC_RELAXED 0 INT_FAST8_MAX __MLIBC_INT_FAST8_MAX INT_FAST16_MAX __MLIBC_INT_FAST16_MAX __has_include_next(STR) __has_include_next__(STR) __VERSION__ "8.2.0" __buffer_ptr __FLT32X_HAS_INFINITY__ 1 __FLT128_HAS_INFINITY__ 1 __MLIBC_INT32_C(x) __INT32_C(x) __UINT_LEAST8_TYPE__ unsigned char __SIZEOF_INT128__ 16 __MLIBC_UINT32_C(x) __UINT32_C(x) __MLIBC_INT_FAST8_MAX __MLIBC_INT8_MAX __MLIBC_CHECK_TYPE(T1,T2) __MLIBC_STATIC_ASSERT(sizeof(T1) == sizeof(T2), #T1 " != " #T2); __INT8_C(c) c PRIiFAST64 "li" __FLT128_MAX__ 1.18973149535723176508575932662800702e+4932F128 ULLONG_MAX (__LONG_LONG_MAX__ * 2ULL + 1ULL) __INT_LEAST32_TYPE__ int __INT_LEAST16_WIDTH__ 16 PRIXLEAST16 "X" UINT64_MAX __MLIBC_UINT64_MAX _T_SIZE_  _GCC_WRAP_STDINT_H  PRIdPTR "ld" _MLIBC_STDINT_H  PRIoLEAST8 "o" ULONG_MAX stdout __unix__ 1 __GCC_HAVE_SYNC_COMPARE_AND_SWAP_1 1 __io_offset __FLT64X_MIN_EXP__ (-16381) __SIZEOF_INT__ 4 _BSD_SIZE_T_  __FLT_DIG__ 6 __INT_FAST16_WIDTH__ 64 WCHAR_MAX __MLIBC_WCHAR_MAX PRIx32 "x" __LDBL_HAS_DENORM__ 1 __MLIBC_UINT_FAST16_C(x) __MLIBC_UINT64_C(x) __DEC32_MIN__ 1E-95DF _POSIX_ARG_MAX 4096 CHAR_BIT 8 __MLIBC_UINT64_C(x) __UINT64_C(x) __GCC_IEC_559 2 __FLT128_MIN_EXP__ (-16381) __FLT32_HAS_QUIET_NAN__ 1 _BSD_SIZE_T_DEFINED_  __UINT_LEAST16_MAX__ 0xffff __UINT_FAST64_MAX__ 0xffffffffffffffffUL PRIXLEAST8 "X" PRIdFAST32 "ld" __UINT_LEAST8_MAX__ 0xff __DEC128_MIN_EXP__ (-6142) INT32_MIN __MLIBC_INT32_MIN __WCHAR_TYPE__ int __INT8_MAX__ 0x7f __GCC_HAVE_SYNC_COMPARE_AND_SWAP_4 1 __need_NULL INT_FAST64_MIN __MLIBC_INT_FAST64_MIN __FLT128_MAX_EXP__ 16384 UINTMAX_MAX __MLIBC_UINTMAX_MAX __FLT_RADIX__ 2 __FLT32X_DENORM_MIN__ 4.94065645841246544176568792868221372e-324F32x UINT_FAST64_MAX __MLIBC_UINT_FAST64_MAX INT_FAST32_MIN __MLIBC_INT_FAST32_MIN __SIZEOF_LONG_DOUBLE__ 16 __DBL_HAS_QUIET_NAN__ 1 INT_LEAST8_MIN __MLIBC_INT8_MIN __MLIBC_UINT8_MAX __UINT8_MAX__ __LDBL_DENORM_MIN__ 3.64519953188247460252840593361941982e-4951L INTMAX_MAX __MLIBC_INTMAX_MAX __FLT64_HAS_INFINITY__ 1 __UINT_FAST8_MAX__ 0xff __ATOMIC_HLE_RELEASE 131072 __LDBL_MAX_EXP__ 16384 __INTMAX_TYPE__ long int MLIBC_SIZE_T_H  INT16_MIN __MLIBC_INT16_MIN __INTPTR_TYPE__ long int __DEC64_MAX__ 9.999999999999999E384DD __MLIBC_INT64_MIN (-__MLIBC_INT64_MAX - 1) __GCC_ATOMIC_INT_LOCK_FREE 2 __MLIBC_UINT_FAST32_C(x) __MLIBC_UINT64_C(x) __MMX__ 1 CHAR_MAX SCHAR_MAX PRIXFAST32 "lX" __FLT64X_DIG__ 18 UINT_LEAST64_MAX __MLIBC_UINT64_MAX __INT_LEAST64_WIDTH__ 64 PRIdFAST64 "ld" __FLT64_MAX_10_EXP__ 308 __ORDER_LITTLE_ENDIAN__ 1234 SHRT_MIN __SIZEOF_PTRDIFF_T__ 8 __DEC128_MANT_DIG__ 34 PRIXPTR "lX" __INT32_TYPE__ int __code_model_small__ 1 __MLIBC_UINT8_C(x) __UINT8_C(x) __FLT64X_HAS_DENORM__ 1 __DEC32_MAX_EXP__ 97 BUFSIZ 512 _IONBF 3 LLONG_MIN (-__LONG_LONG_MAX__ - 1LL) PRIXFAST16 "lX" PRIiLEAST16 "i" __MLIBC_INTPTR_MAX __INTPTR_MAX__ PRIXFAST64 "lX" PRIo16 "o" __MLIBC_INT_FAST64_C(x) __MLIBC_INT64_C(x) __FLT64X_MIN_10_EXP__ (-4931) __MLIBC_UINT_FAST32_MAX __MLIBC_UINT64_MAX __FLT128_MAX_10_EXP__ 4932 __FLT128_MIN__ 3.36210314311209350626267781732175260e-4932F128 PATH_SEPARATOR ':' stdin __FLT64_MIN_10_EXP__ (-307) UINT32_MAX __MLIBC_UINT32_MAX dg_Create __DBL_MAX__ ((double)1.79769313486231570814527423731704357e+308L) __amd64__ 1 PRId16 "d" PRIi64 "li" LLONG_MIN (-LLONG_MAX - 1LL) __FLT32_DECIMAL_DIG__ 9 __FLT128_DIG__ 33 myargc WINT_MAX __MLIBC_WINT_MAX PRIiPTR "li" __WCHAR_WIDTH__ 32 __FLT32_HAS_INFINITY__ 1 __MLIBC_INTMAX_MAX __INTMAX_MAX__ __MLIBC_UINT_FAST64_C(x) __MLIBC_UINT64_C(x) SIG_ATOMIC_MAX __MLIBC_SIG_ATOMIC_MAX __LONG_LONG_MAX__ 0x7fffffffffffffffLL M_FindResponseFile __UINT_LEAST16_TYPE__ short unsigned int __FLT_MAX_10_EXP__ 38 NAME_MAX 255 __LDBL_HAS_INFINITY__ 1 __FLT32X_EPSILON__ 2.22044604925031308084726333618164062e-16F32x NULL ((void *)0) myargv __MLIBC_PTRDIFF_MIN (-__PTRDIFF_MAX__ - 1) PRIi8 "i" _SIZE_T_DEFINED  __INTMAX_MAX__ 0x7fffffffffffffffL D_DoomMain __MLIBC_INT16_C(x) __INT16_C(x) PRIdFAST16 "ld" __FLT64_DECIMAL_DIG__ 17 __SIZEOF_FLOAT128__ 16 __FLT32_MIN_EXP__ (-125) __SIZE_TYPE__ long unsigned int __MLIBC_UINTPTR_MAX __UINTPTR_MAX__ SIZE_MAX __MLIBC_SIZE_MAX __DEC_EVAL_METHOD__ 2 __FLT_MAX__ 3.40282346638528859811704183484516925e+38F __DBL_MIN_10_EXP__ (-307) __MLIBC_INT_FAST16_MAX __MLIBC_INT64_MAX __GXX_ABI_VERSION 1013 __LDBL_MIN_10_EXP__ (-4931) __FLT32_DIG__ 6 __FLT64_HAS_DENORM__ 1 __FLT_EVAL_METHOD__ 0 PRIxFAST64 "lx" ULONG_LONG_MAX __FLT32X_HAS_DENORM__ 1 __x86_64__ 1 __MLIBC_INT_FAST32_MIN __MLIBC_INT64_MIN __INTMAX_C(c) c ## L PTRDIFF_MIN __MLIBC_PTRDIFF_MIN __FLT64X_MAX__ 1.18973149535723176502126385303097021e+4932F64x __DEC64_MIN_EXP__ (-382) __MLIBC_POSIX_OPTION __has_include(<unistd.h>) UCHAR_MAX __SIZE_T__  TMP_MAX 1024 PRIoLEAST16 "o" __INT_LEAST64_MAX__ 0x7fffffffffffffffL __INT_LEAST8_WIDTH__ 8 __UINT8_MAX__ 0xff __UINT16_MAX__ 0xffff LONG_MIN (-LONG_MAX - 1L) _SIZET_  __MLIBC_INT8_C(x) __INT8_C(x) __MLIBC_WINT_MAX __WINT_MAX__ __INT_FAST64_TYPE__ long int __builtin_puts PRIoFAST8 "o" __UINT32_MAX__ 0xffffffffU __INTMAX_WIDTH__ 64 __DEC32_MAX__ 9.999999E96DF UINT_LEAST8_MAX __MLIBC_UINT8_MAX INT32_MAX __MLIBC_INT32_MAX __PTRDIFF_MAX__ 0x7fffffffffffffffL UINT32_C(x) __MLIBC_UINT32_C(x) __INT_LEAST16_TYPE__ short int __FLT32_MAX_EXP__ 128 _BITS_FEATURE_H  PRIuFAST8 "u" UINT16_C(x) __MLIBC_UINT16_C(x) INT_FAST8_MIN __MLIBC_INT_FAST8_MIN __DBL_DIG__ 15 PRIuLEAST64 "lu" __INT_LEAST8_MAX__ 0x7f LLONG_MIN __MLIBC_INT8_MAX __INT8_MAX__ __LP64__ 1 INT32_C(x) __MLIBC_INT32_C(x) LONG_LONG_MIN (-LONG_LONG_MAX - 1LL) __GCC_ATOMIC_LONG_LOCK_FREE 2 __FLT32X_DIG__ 15 __MLIBC_SIG_ATOMIC_MIN __SIG_ATOMIC_MIN__ PRIi32 "i" __FLT32X_MANT_DIG__ 53 PRIdMAX "ld" _ABIBITS_SEEK_WHENCE_H  _LP64 1 INT_MAX __INT_MAX__ __UINT16_TYPE__ short unsigned int __FLT64X_MAX_10_EXP__ 4932 INT16_MAX __MLIBC_INT16_MAX __DBL_MIN__ ((double)2.22507385850720138309023271733240406e-308L) __GCC_ATOMIC_BOOL_LOCK_FREE 2 __UINT_FAST32_MAX__ 0xffffffffffffffffUL __FINITE_MATH_ONLY__ 0 LEMON 1 UCHAR_MAX (SCHAR_MAX * 2 + 1) PRIo8 "o" __MLIBC_STATIC_ASSERT(c,text) _Static_assert(c, text) __FLT64_MAX__ 1.79769313486231570814527423731704357e+308F64 __size_t__  PRIxLEAST8 "x" INT_MIN (-INT_MAX - 1) __MLIBC_ANSI_OPTION __has_include(<stdlib.h>) INT_LEAST64_MAX __MLIBC_INT64_MAX __GCC_ASM_FLAG_OUTPUTS__ 1 __UINT_LEAST64_MAX__ 0xffffffffffffffffUL GNU C17 8.2.0 -mtune=generic -march=x86-64 -ggdb3 -g -Os P_tmpdir "/tmp" PRIu8 "u" __MLIBC_SIZE_MAX __SIZE_MAX__ __ELF__ 1 __FLT32X_MIN__ 2.22507385850720138309023271733240406e-308F32x __UINTPTR_TYPE__ long unsigned int __INT16_C(c) c __GCC_HAVE_DWARF2_CFI_ASM 1 __SIZEOF_FLOAT__ 4 __DEC32_SUBNORMAL_MIN__ 0.000001E-95DF __FLT64X_HAS_QUIET_NAN__ 1 __FLT_HAS_INFINITY__ 1 ULONG_LONG_MAX (LONG_LONG_MAX * 2ULL + 1ULL) PRIXLEAST64 "lX" PRIuLEAST8 "u" PRIx16 "x" _GCC_LIMITS_H_  __STDC__ 1 __SSE2__ 1 PRIo32 "o" INT64_MIN __MLIBC_INT64_MIN __DBL_MAX_EXP__ 1024 __SIZEOF_LONG__ 8 __ATOMIC_CONSUME 1 INT64_MAX __MLIBC_INT64_MAX __USER_LABEL_PREFIX__  __WINT_TYPE__ unsigned int PRIi16 "i" __INT16_MAX__ 0x7fff PRIxFAST32 "lx" __SCHAR_WIDTH__ 8 __UINT32_C(c) c ## U __INT_FAST32_TYPE__ long int PRIxLEAST16 "x" __SIZEOF_DOUBLE__ 8 __GNUC_PATCHLEVEL__ 0 __UINT8_C(c) c __MLIBC_INT16_MAX __INT16_MAX__ __MLIBC_EOF_BIT 1 __WINT_MIN__ 0U PRIoLEAST64 "lo" __LDBL_MANT_DIG__ 64 SEEK_SET 0 __STDC_UTF_16__ 1 __LDBL_EPSILON__ 1.08420217248550443400745280086994171e-19L PRIdLEAST8 "d" PRIuMAX "lu" DIR_SEPARATOR '/' PRIuFAST16 "lu" _GCC_NEXT_LIMITS_H  __INT_FAST8_TYPE__ signed char INT16_C(x) __MLIBC_INT16_C(x) SHRT_MIN (-SHRT_MAX - 1) __GCC_IEC_559_COMPLEX 2 __SIG_ATOMIC_MIN__ (-__SIG_ATOMIC_MAX__ - 1) __MLIBC_INT_FAST64_MIN __MLIBC_INT64_MIN _LIMITS_H___  PRIuPTR "lu" __SIZEOF_WCHAR_T__ 4 PIPE_BUF 4096 __FLT128_MIN_10_EXP__ (-4931) __FLOAT_WORD_ORDER__ __ORDER_LITTLE_ENDIAN__ __GCC_HAVE_SYNC_COMPARE_AND_SWAP_2 1 __DEC32_MANT_DIG__ 7 PRIuFAST32 "lu" __FLT32_DENORM_MIN__ 1.40129846432481707092372958328991613e-45F32 __need_size_t __UINT_FAST16_MAX__ 0xffffffffffffffffUL ULLONG_MAX (LLONG_MAX * 2ULL + 1ULL) __need___va_list __INT32_MAX__ 0x7fffffff ___int_size_t_h  __ATOMIC_ACQUIRE 2 __UINT16_C(c) c LONG_LONG_MAX __LONG_LONG_MAX__ __INT64_MAX__ 0x7fffffffffffffffL __need_size_t  /mnt/e/OneDrive/LemonDOOM/lemondoom PRIoFAST16 "lo" __SEG_GS 1 PRIX32 "X" __SSE_MATH__ 1 CHAR_BIT __UINTMAX_TYPE__ long unsigned int MLIBC_NULL_H  __DEC128_MAX_EXP__ 6145 __MLIBC_INT_FAST32_MAX __MLIBC_INT64_MAX PRIuLEAST16 "u" __SIG_ATOMIC_WIDTH__ 32 __MLIBC_INT_FAST8_MIN __MLIBC_INT8_MIN PRIxMAX "lx" __MLIBC_UINT16_MAX __UINT16_MAX__ __SHRT_MAX__ 0x7fff __GCC_ATOMIC_WCHAR_T_LOCK_FREE 2 UINT_MAX (INT_MAX * 2U + 1U) __ORDER_PDP_ENDIAN__ 3412 UINT8_C(x) __MLIBC_UINT8_C(x) UINT_MAX __MLIBC_UINT_FAST64_MAX __MLIBC_UINT64_MAX PRIxFAST16 "lx" __FLT_DECIMAL_DIG__ 9 PRIxPTR "lx" PRIoFAST64 "lo" __MLIBC_UINT16_C(x) __UINT16_C(x) __LDBL_MIN_EXP__ (-16381) __WINT_WIDTH__ 32 __DEC128_EPSILON__ 1E-33DL __FLT64X_MIN__ 3.36210314311209350626267781732175260e-4932F64x UINT_LEAST16_MAX __MLIBC_UINT16_MAX arrlen(array) (sizeof(array) / sizeof(*array)) __INT_FAST8_MAX__ 0x7f __dirty_end __FLT32_EPSILON__ 1.19209289550781250000000000000000000e-7F32 __x86_64 1 UINT_FAST32_MAX __MLIBC_UINT_FAST32_MAX __LONG_MAX__ 0x7fffffffffffffffL __FLT128_HAS_QUIET_NAN__ 1 __DEC64_MAX_EXP__ 385 PRIu32 "u" INT_LEAST64_MIN __MLIBC_INT64_MIN PRIX64 "lX" __FLT32X_MIN_10_EXP__ (-307) PRId8 "d" PRIdFAST8 "d" __UINTMAX_C(c) c ## UL __DEC64_SUBNORMAL_MIN__ 0.000000000000001E-383DD __MLIBC_INT32_MAX __INT32_MAX__ ULONG_MAX (LONG_MAX * 2UL + 1UL) __FLT64X_HAS_INFINITY__ 1 __DEC128_MIN__ 1E-6143DL __FLT32X_MIN_EXP__ (-1021) __INTPTR_WIDTH__ 64 LONG_BIT (CHAR_BIT * sizeof(long)) __MLIBC_WCHAR_MAX __WCHAR_MAX__ _STRINGS_H  CHAR_MIN SCHAR_MIN __UINT_FAST8_TYPE__ unsigned char __INT32_C(c) c PRIxLEAST64 "lx" __LDBL_HAS_QUIET_NAN__ 1 __INT8_TYPE__ signed char __WINT_MAX__ 0xffffffffU INT8_MIN __MLIBC_INT8_MIN PRIiFAST16 "li" PRIX8 "X" L_tmpnam 256 __UINT32_TYPE__ unsigned int __MLIBC_WCHAR_MIN __WCHAR_MIN__ INT_FAST32_MAX __MLIBC_INT_FAST32_MAX __mlibc_file_base __FLT128_EPSILON__ 1.92592994438723585305597794258492732e-34F128 SCHAR_MIN (-SCHAR_MAX - 1) __offset __SIZEOF_LONG_LONG__ 8 __UINT8_TYPE__ unsigned char __SHRT_WIDTH__ 16 __SSE2_MATH__ 1 PTRDIFF_MAX __MLIBC_PTRDIFF_MAX _T_SIZE  PATH_MAX 4096 UINT_LEAST32_MAX __MLIBC_UINT32_MAX __INT_FAST32_WIDTH__ 64 DIR_SEPARATOR_S "/" _MLIBC_INTERNAL_TYPES_H  PRIxFAST8 "x" PRIx64 "lx" __SIZEOF_POINTER__ 8 __FLT64_EPSILON__ 2.22044604925031308084726333618164062e-16F64 __MLIBC_UINT_FAST16_MIN __MLIBC_UINT64_MIN PRIdLEAST32 "d" __FLT64X_MANT_DIG__ 64 __GNUC_VA_LIST  __WCHAR_MAX__ 0x7fffffff __need___va_list  __FLT_MANT_DIG__ 24 PRIX16 "X" __INT_WIDTH__ 32 __LDBL_DECIMAL_DIG__ 21 __GCC_ATOMIC_POINTER_LOCK_FREE 2 __MLIBC_UINT_FAST64_MIN __MLIBC_UINT64_MIN __SEG_FS 1 __UINT_FAST16_TYPE__ long unsigned int __STDC_VERSION__ 201710L PRIoLEAST32 "o" INT8_C(x) __MLIBC_INT8_C(x) __GCC_ATOMIC_CHAR32_T_LOCK_FREE 2 PRIoFAST32 "lo" ULLONG_MAX __CHAR_BIT__ 8 __valid_limit __ATOMIC_HLE_ACQUIRE 65536 __STDC_HOSTED__ 1 PRId64 "ld" __SIZE_WIDTH__ 64 LLONG_MAX __LONG_LONG_MAX__ __has_include(STR) __has_include__(STR) __MLIBC_INT_FAST64_MAX __MLIBC_INT64_MAX MLIBC_OFF_T_H  INTMAX_MIN __MLIBC_INTMAX_MIN __LONG_WIDTH__ 64 __UINT64_MAX__ 0xffffffffffffffffUL INT_LEAST8_MAX __MLIBC_INT8_MAX PRIu16 "u" LONG_MAX __LONG_MAX__ __k8 1 __GCC_ATOMIC_LLONG_LOCK_FREE 2 __FLT_MAX_EXP__ 128 __ATOMIC_ACQ_REL 4 MLIBC_SSIZE_T_H  __MLIBC_UINT_FAST16_MAX __MLIBC_UINT64_MAX __DEC32_MIN_EXP__ (-94) PRIu64 "lu" __INT64_TYPE__ long int __FLT_MIN__ 1.17549435082228750796873653722224568e-38F INTPTR_MAX __MLIBC_INTPTR_MAX PRIoMAX "lo" INT_FAST16_MIN __MLIBC_INT_FAST16_MIN __MLIBC_WINT_MIN __WINT_MIN__ __MLIBC_PTRDIFF_MAX __PTRDIFF_MAX__ __FXSR__ 1 PRIoPTR "lo" __INT_LEAST32_WIDTH__ 32 UINT_FAST16_MAX __MLIBC_UINT_FAST16_MAX __UINTMAX_MAX__ 0xffffffffffffffffUL INT_LEAST32_MIN __MLIBC_INT32_MIN PRIiLEAST8 "i" INT_LEAST16_MAX __MLIBC_INT16_MAX UINT_FAST8_MAX __MLIBC_UINT_FAST8_MAX __MLIBC_ERROR_BIT 2 CHAR_BIT __CHAR_BIT__ __MLIBC_UINT_FAST32_MIN __MLIBC_UINT64_MIN __UINT_LEAST64_TYPE__ long unsigned int __lemon__ 1 PRIXLEAST32 "X" __MLIBC_INT16_MIN (-__MLIBC_INT16_MAX - 1) __status_bits __MLIBC_UINT_FAST8_C(x) __MLIBC_UINT8_C(x) __SIZE_MAX__ 0xffffffffffffffffUL PACKEDATTR __attribute__((packed)) __GCC_ATOMIC_SHORT_LOCK_FREE 2 __FLT64X_DECIMAL_DIG__ 21 __OPTIMIZE_SIZE__ 1 __INT_FAST16_MAX__ 0x7fffffffffffffffL NORMALUNIX 1 __FLT_EPSILON__ 1.19209289550781250000000000000000000e-7F __FLT_EVAL_METHOD_TS_18661_3__ 0 __DBL_HAS_INFINITY__ 1 INT_LEAST16_MIN __MLIBC_INT16_MIN __INT64_C(c) c ## L __MLIBC_UINT_FAST8_MIN __MLIBC_UINT8_MIN __MLIBC_INT_FAST16_C(x) __MLIBC_INT64_C(x) INT_FAST64_MAX __MLIBC_INT_FAST64_MAX SCHAR_MAX __SCHAR_MAX__ __FLT64_MIN_EXP__ (-1021) __PTRDIFF_TYPE__ long int __DOOMTYPE__  __INT_FAST16_TYPE__ long int PRIo64 "lo" __DEC128_SUBNORMAL_MIN__ 0.000000000000000000000000000000001E-6143DL __MLIBC_UINT32_MAX __UINT32_MAX__ __MLIBC_UINTMAX_MAX __UINTMAX_MAX__ MB_LEN_MAX 1 PRIiFAST8 "i" _SIZE_T_DECLARED  __SIZEOF_FLOAT80__ 16 __FLT32X_HAS_QUIET_NAN__ 1 __DBL_MAX_10_EXP__ 308 __GCC_ATOMIC_CHAR_LOCK_FREE 2 __GNUC_STDC_INLINE__ 1 __SSE__ 1 __MLIBC_INT64_MAX __INT64_MAX__ __BIGGEST_ALIGNMENT__ 16 __FLT128_DENORM_MIN__ 6.47517511943802511092443895822764655e-4966F128 _SYS_SIZE_T_H  __MLIBC_INTPTR_MIN (-__INTPTR_MAX__ - 1) __MLIBC_INT_FAST8_C(x) __MLIBC_INT8_C(x) PRIdLEAST64 "ld" __FLT_MIN_EXP__ (-125) UINT16_MAX __MLIBC_UINT16_MAX SCNu64 "lu" __size_t  __DEC128_MAX__ 9.999999999999999999999999999999999E6144DL __REGISTER_PREFIX__  USHRT_MAX LONG_LONG_MIN PRIuLEAST32 "u" __UINT_LEAST32_MAX__ 0xffffffffU __FLT32X_MAX_10_EXP__ 308 __amd64 1 __M_ARGV__  LINE_MAX 4096 UINTPTR_MAX __MLIBC_UINTPTR_MAX __MLIBC_UINT64_MAX __UINT64_MAX__ __FLT64_DENORM_MIN__ 4.94065645841246544176568792868221372e-324F64 __FLT32_MAX_10_EXP__ 38 __dirty_begin __FLT128_DECIMAL_DIG__ 36 __PTRDIFF_WIDTH__ 64 __INT_LEAST32_MAX__ 0x7fffffff SHRT_MAX __SHRT_MAX__ __UINT_FAST64_TYPE__ long unsigned int PRIx8 "x" __LDBL_MAX_10_EXP__ 4932 __DEC64_MIN__ 1E-383DD __FLT32_MIN__ 1.17549435082228750796873653722224568e-38F32 __DBL_EPSILON__ ((double)2.22044604925031308084726333618164062e-16L) PRIiLEAST64 "li" __PRAGMA_REDEFINE_EXTNAME 1 __SIG_ATOMIC_TYPE__ int __FLT64X_DENORM_MIN__ 3.64519953188247460252840593361941982e-4951F64x PRId32 "d" __FLT128_HAS_DENORM__ 1 USHRT_MAX (SHRT_MAX * 2 + 1) INT64_C(x) __MLIBC_INT64_C(x) __INT_FAST8_WIDTH__ 8 __MLIBC_LINUX_OPTION __has_include(<linux/types.h>) __FLT64_MANT_DIG__ 53 __DEC64_MANT_DIG__ 16 __FLT_HAS_DENORM__ 1 __INT_FAST64_WIDTH__ 64 __DECIMAL_DIG__ 21 dummy.c net_client_connected drone true I_InitTimidityConfig boolean false undef ssecret totalitems THUSTR_7 "level 7: prison" C3TEXT "YOU ARE AT THE CORRUPT HEART OF THE CITY,\n""SURROUNDED BY THE CORPSES OF YOUR ENEMIES.\n""YOU SEE NO WAY TO DESTROY THE CREATURES'\n""ENTRYWAY ON THIS SIDE, SO YOU CLENCH YOUR\n""TEETH AND PLUNGE THROUGH IT.\n""\n""THERE MUST BE A WAY TO CLOSE IT ON THE\n""OTHER SIDE. WHAT DO YOU CARE IF YOU'VE\n""GOT TO GO THROUGH HELL TO GET TO IT?" SPR_LAUN exe_final2 SPR_PUNG S_BOS2_RAISE1 S_BOS2_RAISE2 S_BOS2_RAISE3 S_BOS2_RAISE4 S_BOS2_RAISE5 S_BOS2_RAISE6 S_BOS2_RAISE7 WALLRANGE REDRANGE maxkills momx momy momz GRAYSRANGE 16 KEY_EQUALS 0x3d MAXSPECIALCROSS_ORIGINAL 8 CC_ZOMBIE "ZOMBIEMAN" evtype_t CC_HELL "HELL KNIGHT" HUSTR_TALKTOSELF5 "You've lost it..." CDWALLRANGE YELLOWRANGE waiting SPR_MGUN S_SKEL_PAIN levelTimer S_VILE_DIE2 data1 data2 S_FATT_RUN3 data4 S_VILE_DIE8 MT_TRACER S_FATT_RUN8 S_BRAINEYE1 S_BSPI_STND HUSTR_28 "level 28: the spirit world" middle AM_changeWindowScale S_PINS2 S_DSNR1 S_PINS4 S_HANGTSKULL centerxfrac GOTBLUESKUL "Picked up a blue skull key." S_DSGUN10 S_ARM1A MAXBUTTONS 16 THUSTR_26 "level 26: ballistyx" PU_SOUND AM_clipMline S_PVIS MAXRADIUS 32*FRACUNIT NET_RELIABLE_PACKET (1 << 15) bnext S_PLASMADOWN __V_VIDEO__  ANG1 (ANG45 / 45) blazeDWUS T1TEXT "You've fought your way out of the infested\n""experimental labs.   It seems that UAC has\n""once again gulped it down.  With their\n""high turnover, it must be hard for poor\n""old UAC to buy corporate health insurance\n""nowadays..\n""\n""Ahead lies the military complex, now\n""swarming with diseased horrors hot to get\n""their teeth into you. With luck, the\n""complex still has some warlike ordnance\n""laying around." S_PMAP S_MISSILE S_SAWB GOTINVIS "Partial Invisibility" AM_restoreScaleAndLoc S_PLASMA1 S_PLASMA2 sfxVolume viewangleoffset S_SARG_RUN1 S_SARG_RUN2 S_ARM2A iquehead S_SARG_RUN5 S_SARG_RUN6 S_SARG_RUN7 S_SARG_RUN8 soundorg fullscreen va_end(v) __builtin_va_end(v) key_menu_quit S_MISSILEUP midtexture sscount VDOORWAIT 150 QSAVESPOT "you haven't picked a quicksave slot yet!\n\n"PRESSKEY S_TROO_STND mousebjump textureheight T3TEXT "The vista opening ahead looks real damn\n""familiar. Smells familiar, too -- like\n""fried excrement. You didn't like this\n""place before, and you sure as hell ain't\n""planning to like it now. The more you\n""brood on it, the madder you get.\n""Hefting your gun, an evil grin trickles\n""onto your face. Time to take some names." HUSTR_E1M5 "E1M5: Phobos Lab" WHITE (256-47) PHUSTR_11 "level 11: hunted" MTF_EASY 1 S_CPOS_RAISE1 S_CPOS_RAISE2 S_CPOS_RAISE3 key_useartifact S_CPOS_RAISE5 S_CPOS_RAISE6 S_CPOS_RAISE7 S_SKULL_DIE5 S_SKULL_DIE6 sprev __I_SYSTEM__  HUSTR_TALKTOSELF1 "You mumble to yourself" readyweapon bottomtexture S_RSKULL soundtraversed AM_clearFB S_GTORCHSHRT2 S_GTORCHSHRT3 S_GTORCHSHRT4 S_BTORCHSHRT key_message_refresh spawnstate stime CC_SHOTGUN "SHOTGUN GUY" wp_bfg S_BSKULL HUSTR_25 "level 25: bloodfalls" DEH_VANILLA_NUMSFX 107 STSTR_KFAADDED "Very Happy Ammo Added" SPR_SAWG PHUSTR_18 "level 18: neurosphere" PU_FREE lastspritelump S_BSPI_ATK1 S_BSPI_ATK2 S_BSPI_ATK3 AM_Start key_menu_up S_PAIN_DIE1 S_PAIN_DIE2 S_PAIN_DIE3 S_PAIN_DIE4 S_PAIN_DIE5 S_PAIN_DIE6 mousebforward SPR_GOR1 SPR_GOR2 SPR_GOR3 SPR_GOR4 SPR_GOR5 S_BRAIN_PAIN drawsegs S_MISSILEFLASH1 BLUES (256-4*16+8) S_MISSILEFLASH3 S_SGUN damagecount SPR_CBRA S_PVIS2 THUSTR_8 "level 8: metal" pw_invulnerability KEYP_7 KEY_HOME S_CYBER_PAIN S_KEENPAIN2 colormaps S_SPID_ATK2 S_SPID_ATK3 S_NULL MT_SHADOWS GAMMALVL3 "Gamma correction level 3" TSWALLCOLORS GRAYS KEY_F8 (0x80+0x42) key_strafe HUSTR_CHATMACRO3 "I'm not looking too good!" D_CDROM "CD-ROM Version: default.cfg from c:\\doomdata\n" NET_DEFS_H  S_PLASMA extralight MT_POSSESSED finit_height MAPBMASK (MAPBLOCKSIZE-1) S_BRAINEYESEE consoleplayer PHUSTR_14 "level 14: genesis" S_BOSS_RAISE1 S_BOSS_RAISE2 S_BOSS_RAISE3 S_BOSS_RAISE4 S_BOSS_RAISE5 S_BOSS_RAISE6 S_BOSS_RAISE7 lumpinfo_s lumpinfo_t S_TROO_ATK1 S_TROO_ATK2 S_TROO_ATK3 upstate __P_MOBJ__  MAX_DM_STARTS 10 GOTINVUL "Invulnerability!" key_menu_help in_stasis THUSTR_6 "level 6: open season" LIGHTSEGSHIFT 4 PHUSTR_31 "level 31: cyberden" plat_e CC_SPIDER "THE SPIDER MASTERMIND" NUMWEAPONS S_ARM1 S_ARM2 fastCrushAndRaise viewplayer arti HUSTR_MESSAGESENT "[Message Sent]" intercept_p key_arti_all S_STIM key_menu_right SPR_BROK key_menu_load KEY_DOWNARROW 0xaf S_SPOS_XDIE1 S_SPOS_XDIE2 S_SPOS_XDIE3 S_SPOS_XDIE4 S_SPOS_XDIE5 S_SPOS_XDIE6 S_SPOS_XDIE7 S_SPOS_XDIE8 S_SPOS_XDIE9 event_t SPR_KEEN S_DEADTORSO SPR_MISF SPR_MISG SPR_MISL blockmaplump key_flyup demoplayback KEYP_2 KEY_DOWNARROW HUSTR_E1M9 "E1M9: Military Base" PHUSTR_27 "level 27: anti-christ" MAXPLATS 30 T5TEXT "What now? Looks totally different. Kind\n""of like King Tut's condo. Well,\n""whatever's here can't be any worse\n""than usual. Can it?  Or maybe it's best\n""to let sleeping gods lie.." finit_width MTOF(x) (FixedMul((x),scale_mtof)>>16) GOTSUIT "Radiation Shielding Suit" key_menu_decscreen weaponowned cards m_paninc EMPTYSTRING "empty slot" AM_drawGrid sidenum KEY_F2 (0x80+0x3c) bottomheight ds_colormap joybstrafe S_SAW pw_allmap QLOADNET "you can't quickload during a netgame!\n\n"PRESSKEY frontsector PHUSTR_30 "level 30: the gateway of hell" S_MEAT2 S_MEAT3 S_MEAT4 joybnextweapon GameMode_t S_PLASMAUP REDRANGE 16 S_PISTOL S_EVILEYE NUMSPRITES HUSTR_E2M3 "E2M3: Refinery" S_PLAY_ATK1 S_PLAY_ATK2 rw_angle1 bmaporgx bmaporgy yslope am_misl S_BEXP2 S_BEXP3 S_BEXP4 ceiling_e floorfunc S_STALAGTITE SPR_BRS1 R (FRACUNIT) think_t doomednum CC_BARON "BARON OF HELL" AM_loadPics E2TEXT "You've done it! The hideous cyber-\n""demon lord that ruled the lost Deimos\n""moon base has been slain and you\n""are triumphant! But ... where are\n""you? You clamber to the edge of the\n""moon and look down to see the awful\n""truth.\n" "\n""Deimos floats above Hell itself!\n""You've never heard of anyone escaping\n""from Hell, but you'll make the bastards\n""sorry they ever heard of you! Quickly,\n""you rappel down to  the surface of\n""Hell.\n""\n" "Now, it's on to the final chapter of\n""DOOM! -- Inferno." am_map.c armorpoints NIGHTMARE "are you sure? this skill level\n""isn't even remotely fair.\n\n"PRESSYN scale_ftom S_SGUNDOWN VDOORSPEED FRACUNIT*2 HUSTR_CHATMACRO8 "I'll take care of it." GOTREDSKULL "Picked up a red skull key." HUSTR_KEYBROWN 'b' MT_MISC7 MT_MISC8 MT_MISC9 screenvisible rowoffset finecosine S_PLASBALL lightlev scale1 scale2 key_right gamestate_t DEH_String(x) (x) powers S_BSPI_DIE1 MAXLIGHTSCALE 48 SPR_COL1 SPR_YSKU SPR_COL3 SPR_COL4 SPR_COL5 SPR_COL6 bwhere_e skymap mobj_s S_SHRTGRNCOL data3 THUSTR_27 "level 27: mount pain" HUSTR_24 "level 24: the chasm" SPR_COLU heretic GOTMEDINEED "Picked up a medikit that you REALLY need!" markpoints HUSTR_E3M6 "E3M6: Mt. Erebus" S_VILE_ATK5 STSTR_FAADDED "Ammo (no keys) Added" numsprites states sequence_len maskedtexturecol flashstate wp_fist viewwindowy S_ROCKET deltaviewheight __INFO__  sk_noitems FixedDiv HUSTR_E3M2 "E3M2: Slough of Despair" PHUSTR_25 "level 25: the temple of darkness" dc_yh S_FATSHOTX1 S_FATSHOTX2 dc_yl gamedescription SCREENWIDTH 320 pw_ironfeet HUSTR_E4M2 "E4M2: Perfect Hatred" demorecording GOTCHAINSAW "A chainsaw!  Find some meat!" S_BLOODYTWITCH2 S_PLASMAFLASH1 S_PLASMAFLASH2 __R_THINGS__  FF_FRAMEMASK 0x7fff S_TROO_DIE2 S_TROO_DIE3 S_TROO_DIE4 S_TROO_DIE5 joybspeed HUSTR_E3M3 "E3M3: Pandemonium" HUSTR_TALKTOSELF3 "You scare yourself" lookfly S_SPOS_RUN1 S_SPOS_RUN2 S_SPOS_RUN4 MT_INS S_SPOS_RUN7 MT_INV S_BRAINEYE key_map_mark S_POSS_DIE4 deh_apply_cheats score joybfire S_SPID_STND GREENS (7*16) MAXDRAWSEGS 256 MAX_CHEAT_PARAMS 5 key_invend clipangle MT_BRUISER S_SKEL_DIE5 THUSTR_2 "level 2: human bbq" buttons2 S_VILE_PAIN2 S_COMMKEEN11 S_COMMKEEN12 key_invright S_BON1 armortype S_CPOS_PAIN2 THUSTR_14 "level 14: steel works" SPR_APBX bigstate NUMPOWERS AM_Stop key_menu_forward THUSTR_10 "level 10: redemption" GOTROCKBOX "Picked up a box of rockets." SAVEGAMENAME "doomsav" FEATURE_WAD_MERGE SPR_BKEY HUSTR_E4M3 "E4M3: Sever The Wicked" min_w GOTSUPER "Supercharge!" it_yellowcard AM_rotate M_ZOOMOUT ((int) (FRACUNIT/1.02)) THUSTR_21 "level 21: administration center" player_s S_HEADSONSTICK FixedMul S_BFG1 S_BFG2 S_BFG3 S_BFG4 MT_FIRE S_COLONGIBS leftoffset S_TBALLX1 S_TBALLX2 S_TBALLX3 skills GOTSTIM "Picked up a stimpack." lowfloor KEY_FIRE 0xa3 S_BSPI_ATK4 PT_EARLYOUT 4 S_TFOG S_MISSILE1 S_MISSILE2 S_MISSILE3 AM_Responder fuck FF_FULLBRIGHT 0x8000 S_BOSS_PAIN HUSTR_PLRINDIGO "Indigo: " GOTYELWCARD "Picked up a yellow keycard." STSTR_NOMUS "IMPOSSIBLE SELECTION" savegamedir S_SKEL_MISS1 S_SKEL_MISS2 S_PUNCH WALLCOLORS REDS S_SPID_STND2 refire cheat_player_arrow NET_TICDIFF_SIDE (1 << 1) HUSTR_29 "level 29: the living end" S_FATT_PAIN levelstarttic S_PLAY_DIE1 S_PLAY_DIE2 S_PLAY_DIE3 S_PLAY_DIE4 S_PLAY_DIE5 S_PLAY_DIE6 negonearray oldstatus MT_PAIN MT_MISC11 MT_MISC13 NUMAMMO KEY_LALT KEY_RALT MT_MISC15 wp_plasma centery itemcount their_color floorplane numspritelumps exe_doom_1_2 exe_doom_1_7 exe_doom_1_8 exe_doom_1_9 S_SPID_ATK4 colorrange HUSTR_E2M1 "E2M1: Deimos Anomaly" HUSTR_E2M6 "E2M6: Halls of the Damned" key_invpop atkstate KEYP_5 '5' S_SGUNFLASH1 S_SGUNFLASH2 exe_ultimate psprites key_up S_CLIP gametic key_mission MT_MISC22 GAMMALVL0 "Gamma correction OFF" MT_ARACHPLAZ NUMMOBJTYPES S_SARG_STND vissprite_s vissprite_t S_FATT_PAIN2 S_IFOG01 S_IFOG02 screen_bpp vissprites AM_drawWalls blocklinks lastepisode toptexture SPR_SPOS KEY_RCTRL (0x80+0x1d) S_SPOS_STND S_DSGUN clipammo key_map_north YOURRANGE 0 KEY_F9 (0x80+0x43) THUSTR_18 "level 18: mill" GOTMAP "Computer Area Map" S_TROO_PAIN2 snd_DesiredSfxDevice MAPBLOCKSHIFT (FRACBITS+7) KEY_SCRLCK (0x80+0x46) THUSTR_23 "level 23: lunar mining project" MAXINTERCEPTS (MAXINTERCEPTS_ORIGINAL + 61) ONCEILINGZ INT_MAX S_SPID_DIE5 S_HEAD_RAISE6 SPR_RSKU S_TORCHTREE PLATSPEED FRACUNIT KEY_INS (0x80+0x52) key_straferight MT_MISC10 MT_MISC12 flattranslation MT_MISC14 NET_TICDIFF_FORWARD (1 << 0) MT_MISC16 MT_MISC17 MT_MISC18 MT_MISC19 openrange C6TEXT "CONGRATULATIONS, YOU'VE FOUND THE\n""SUPER SECRET LEVEL!  YOU'D BETTER\n""BLAZE THROUGH THIS ONE!\n" mousebbackward min_scale_mtof CC_REVEN "REVENANT" AMSTR_MARKEDSPOT "Marked Spot" S_BSPI_PAIN2 S_FIRE1 S_FIRE2 S_FIRE4 S_FIRE5 S_FIRE6 S_FIRE7 key_menu_volume S_FIRE9 THUSTR_5 "level 5: hanger" S_PUFF2 it_yellowskull MT_BLOOD movecount HUSTR_E2M4 "E2M4: Deimos Lab" exe_final MT_MISC20 MT_MISC21 __R_PLANE__  MT_MISC23 MT_MISC24 MT_MISC25 MT_MISC26 MT_MISC27 MT_MISC28 MT_MISC29 S_TROO_DIE1 testcontrols_mousespeed outcode1 S_SSWV_RUN1 S_SSWV_RUN2 S_SSWV_RUN3 S_SSWV_RUN5 S_SSWV_RUN6 S_SSWV_RUN7 S_SSWV_RUN8 totalkills FRACUNIT (1<<FRACBITS) wp_pistol PU_LEVEL S_PLAY_XDIE1 S_PLAY_XDIE2 S_PLAY_XDIE3 S_PLAY_XDIE4 S_PLAY_XDIE5 S_PLAY_XDIE6 S_PLAY_XDIE7 S_PLAY_XDIE8 S_PLAY_XDIE9 key_arti_egg ds_xfrac NET_MAGIC_NUMBER 3436803284U FRACBITS 16 GOTBACKPACK "Picked up a backpack full of ammo!" key_flydown sprtopclip MT_MISC30 MT_MISC32 MT_MISC33 MT_MISC34 MT_MISC35 MT_MISC36 mobjtype_t MT_MISC38 MT_MISC39 SPR_CSAW S_SARG_ATK1 S_SARG_ATK2 S_SARG_ATK3 NET_TICDIFF_RAVEN (1 << 6) S_SOUL2 S_SOUL3 S_SOUL4 S_SOUL5 S_SOUL6 key_jump KEYP_MINUS '-' key_menu_back S_BLOOD2 S_HEADCANDLES S_BLOOD3 logical_gamemission (gamemission == pack_chex ? doom : gamemission == pack_hacx ? doom2 : gamemission) painchance MT_MISC40 displayplayer MT_MISC42 MT_MISC43 MT_MISC46 actionf_v MT_MISC49 SPR_APLS SPR_PISF skill_t xtoviewangle KEY_F3 (0x80+0x3d) ev_keydown key_menu_endgame S_BSPI_RAISE1 S_BSPI_RAISE2 S_BSPI_RAISE3 S_BOSS_DIE4 S_BSPI_RAISE5 KEY_RSHIFT (0x80+0x36) S_BSPI_RAISE7 S_SSWV_XDIE5 S_SSWV_XDIE6 S_SSWV_XDIE7 S_SSWV_XDIE8 S_SSWV_XDIE9 KEYP_8 KEY_UPARROW W_ReleaseLumpName KEYP_4 KEY_LEFTARROW MT_BFG MT_MISC50 MT_MISC52 MT_MISC53 MT_MISC54 MT_MISC55 MT_MISC56 MT_MISC57 MT_MISC58 MT_MISC59 S_BKEY2 SPR_BOS2 registered S_BON1C S_BOSS_STND SPR_CHGF SPR_CHGG MT_BARREL S_BEXP5 S_TECHLAMP2 HUSTR_10 "level 10: refueling base" __D_STATE__  S_FATSHOTX3 MT_MISC60 MT_MISC61 AM_initVariables MT_MISC63 MT_MISC64 MT_MISC65 MT_MISC66 MT_MISC67 MT_MISC68 MT_MISC69 MELEERANGE (64*FRACUNIT) snd_MusicDevice SPR_SGN2 raiseToHighest MT_MISC41 MT_SPAWNFIRE Z_ChangeTag(p,t) Z_ChangeTag2((p), (t), __FILE__, __LINE__) SPR_FBXP MT_MISC48 HUSTR_PLRGREEN "Green: " dc_texturemid key_map_maxzoom __mlibc_uint8 S_SBOX MT_MISC70 MT_MISC72 MT_MISC73 MT_MISC74 MT_MISC75 MT_MISC76 MT_BOSSSPIT MT_MISC78 MT_MISC79 PT_ADDLINES 1 THUSTR_29 "level 29: river styx" KEYP_DIVIDE '/' AM_changeWindowLoc S_BON2A S_BON2B key_invleft chatchar S_IFOG MAPBTOFRAC (MAPBLOCKSHIFT-FRACBITS) S_SPID_DIE1 S_SPID_DIE2 S_SPID_DIE3 S_SPID_DIE4 S_SPID_DIE6 S_SPID_DIE7 S_SPID_DIE8 S_SPID_DIE9 max_scale_mtof fline_t PHUSTR_3 "level 3: aztec" playerstarts translationtables secretcount cheat_choppers key_use drawseg_s MT_MISC81 MT_MISC82 MT_MISC83 MT_MISC84 MT_MISC85 MT_MISC86 BROWNS (4*16) MT_HEAD __I_VIDEO__  PHUSTR_2 "level 2: well of souls" GOTMEGA "Picked up the MegaArmor!" MAXCEILINGS 30 numspechit mousebnextweapon mouseSensitivity HUSTR_E4M5 "E4M5: They Will Repent" HUSTR_E1M2 "E1M2: Nuclear Plant" KEY_MINUS 0x2d S_DSGUNDOWN ftom_zoommul S_CYBER_DIE10 S_SARG_STND2 S_PAIN_ATK3 __Z_ZONE__  KEYP_6 KEY_RIGHTARROW HUSTR_E3M8 "E3M8: Dis" ITEMQUESIZE 128 NUM_QUITMESSAGES 8 startmap S_BFUG SPR_PVIS FLOORSPEED FRACUNIT __R_STATE__  min_y SPR_PMAP sprbottomclip subsector_s S_SKEL_PAIN2 THUSTR_31 "level 31: pharaoh" AM_drawLineCharacter S_BSPI_SIGHT downWaitUpStay HUSTR_5 "level 5: the waste tunnels" startfrac flip HUSTR_1 "level 1: entryway" sitems S_FATSHOT1 S_FATSHOT2 PHUSTR_4 "level 4: caged" GOTPLASMA "You got the plasma gun!" finetangent PUTDOT(xx,yy,cc) fb[(yy)*f_w+(xx)]=(cc) gamemap __P_SPEC__  S_STALAG playerstate_t KEY_CAPSLOCK (0x80+0x3a) S_RBALL1 S_RBALL2 STROBEBRIGHT 5 S_HANGBNOBRAIN S_MISSILEDOWN dc_translation SLOPERANGE 2048 key_map_clearmark HUSTR_E1M6 "E1M6: Central Processing" mousebstrafeleft function __W_WAD__  MT_SHOTGUN MT_SHOTGUY CC_HERO "OUR HERO" MT_TROOP S_BOS2_RUN1 S_BOS2_RUN2 S_BOS2_RUN3 S_BOS2_RUN4 S_BOS2_RUN5 S_BOS2_RUN6 S_BOS2_RUN7 S_BOS2_RUN8 MT_MISC62 GS_INTERMISSION islp MO_TELEPORTMAN 14 btexture __M_MISC__  S_SARG_DIE1 S_SARG_DIE2 S_SARG_DIE3 S_SARG_DIE4 S_SARG_DIE5 S_SARG_DIE6 S_POSS_RUN1 S_POSS_RUN2 S_POSS_RUN3 S_POSS_RUN4 S_POSS_RUN5 S_POSS_RUN6 S_POSS_RUN7 S_POSS_RUN8 S_DSGUNUP hscalelight deh_allow_extended_strings S_FATT_RUN7 S_VILE_DIE7 BACKUPTICS 128 S_VILE_DIE9 rw_normalangle it_redcard S_TECHPILLAR KEY_STRAFE_R 0xa1 _STDARG_H  MSGOFF "Messages OFF" ANG1_X 0x01000000 ST_Y (SCREENHEIGHT - ST_HEIGHT) firstline wp_chaingun islope_t m_y2 pack_plut HUSTR_17 "level 17: tenements" spawnpoint actionf_p2 ML_TWOSIDED 4 S_LIVESTICK2 S_SKEL_FIST1 S_SKEL_FIST3 S_SKEL_FIST4 KEY_F11 (0x80+0x57) numlines topheight S_SKULL_STND S_PAIN_PAIN side_t KEY_PRTSCR (0x80+0x59) line_s PD_BLUEO "You need a blue key to activate this object" S_FATT_DIE1 S_FATT_DIE2 ds_yfrac old_m_h strife SCREENHEIGHT 200 S_FATT_DIE5 cht_CheckCheat PU_MUSIC old_m_w old_m_y S_VILE_RUN3 S_VILE_RUN4 S_VILE_RUN5 S_VILE_RUN6 S_VILE_RUN7 S_PMAP4 S_VILE_RUN9 readystate S_BFG MT_MISC77 __D_TICCMD__  S_FATT_RUN12 SPR_TBLU SPR_BBRN S_HEAD_STND S_LIVESTICK dc_iscale AMSTR_GRIDOFF "Grid OFF" THUSTR_1 "level 1: system control" spanfunc S_AMMO FDWALLCOLORS BROWNS THUSTR_20 "level 20: central processing" numframes __D_EVENT__  litelevelscnt SPR_ARM1 SPR_ARM2 SIL_NONE 0 S_VILE_RUN10 S_VILE_RUN11 S_VILE_RUN12 CC_ARCH "ARCH-VILE" S_SARG_RUN4 xiscale S_SPAWNFIRE1 S_SPAWNFIRE3 S_SPAWNFIRE4 S_SPAWNFIRE5 S_SPAWNFIRE6 S_SPAWNFIRE7 scalelightfixed SPR_STIM STSTR_BEHOLDX "Power-up Toggled" THUSTR_30 "level 30: last call" S_SAWUP AM_unloadPics S_BRAIN_DIE1 S_RBALLX1 S_RBALLX2 S_RBALLX3 KEY_DEL (0x80+0x53) usergame automapactive thinker_s inventory MT_BOSSBRAIN ML_DONTPEGTOP 8 STSTR_NCON "No Clipping Mode ON" S_HEAD_DIE4 S_YSKULL nomonsters pspritescale R ((8*PLAYERRADIUS)/7) __DOOMKEYS__  S_BTORCHSHRT3 basecolfunc MT_TROOPSHOT AM_minOutWindowScale AMSTR_FOLLOWON "Follow Mode ON" __va_copy(d,s) __builtin_va_copy(d,s) HUSTR_22 "level 22: the catacombs" S_SPOS_ATK1 S_SPOS_ATK2 S_SPOS_ATK3 S_SKEL_STND2 planefunction_t S_MEGA2 S_MEGA3 S_MEGA4 S_BFGEXP2 S_BFGEXP3 S_BFGEXP4 S_VILE_ATK11 S_SKULL_ATK4 S_BBAR1 S_BBAR2 S_BBAR3 QLPROMPT "do you want to quickload the game named\n\n'%s'?\n\n"PRESSYN mousebprevweapon S_ARACH_PLAZ AM_Ticker _VA_LIST_DEFINED  S_POSS_STND2 S_POSS_RAISE1 S_POSS_RAISE2 S_POSS_RAISE3 S_POSS_RAISE4 S_GIBS __M_FIXED__  lastlook attacker HUSTR_E4M1 "E4M1: Hell Beneath" S_TROO_XDIE5 S_TROO_XDIE6 S_TROO_XDIE7 key_multi_msgplayer key_weapon1 S_HEAD_ATK1 S_HEAD_ATK2 S_HEAD_ATK3 AM_Drawer D_DEVSTR "Development mode ON.\n" raisestate PHUSTR_7 "level 7: caughtyard" ST_Responder S_BLUETORCH2 S_BLUETORCH3 S_BLUETORCH4 SPR_BEXP FINEMASK (FINEANGLES-1) mass PHUSTR_17 "level 17: compound" S_SHRTREDCOL CYMTOF(y) (f_y + (f_h - MTOF((y)-m_y))) S_BOS2_PAIN2 FINEANGLES 8192 SPR_SKEL centerx testcontrols CC_DEMON "DEMON" actionf_p1 S_HEAD_RUN1 S_FATT_RUN10 S_FATT_RUN11 S_CELP key_invdrop SPR_POL3 SPR_POL4 THUSTR_15 "level 15: dead zone" I_VideoBuffer spryscale __TABLES__  GOTROCKET "Picked up a rocket." SPR_POB1 SPR_POB2 KEY_F4 (0x80+0x3e) TICRATE 35 MT_SERGEANT deh_allow_long_cheats S_PLASBALL2 GOTSHOTGUN "You got the shotgun!" S_BRAINSTEM THUSTR_25 "level 25: baron's den" screen_height S_SKEL_MISS3 S_SKEL_MISS4 vsprsortedhead lineguy KEY_END (0x80+0x4f) ML_DONTPEGBOTTOM 16 key_menu_messages S_RKEY pack_hacx sidemove dirtybox S_ARACH_PLEX S_SSWV_STND SPR_SPID S_VILE_HEAL1 S_VILE_HEAL2 PU_LEVSPEC __D_PLAYER__  HUSTR_6 "level 6: the crusher" DEH_MAIN_H  S_VILE_RUN8 wp_supershotgun pad1 S_BSPI_PAIN gameversion pad4 S_FATT_ATK10 HUSTR_CHATMACRO6 "Next time, scumbag..." S_SPID_PAIN2 T2TEXT "You hear the grinding of heavy machinery\n""ahead.  You sure hope they're not stamping\n""out new hellspawn, but you're ready to\n""ream out a whole herd if you have to.\n""They might be planning a blood feast, but\n""you feel about as mean as two thousand\n""maniacs packed into one mad killer.\n""\n""You don't plan to go down easy." it_blueskull S_BSPI_RUN10 S_BSPI_RUN11 S_BSPI_RUN12 activeplats CC_LOST "LOST SOUL" key_menu_qload S_PMAP2 S_PMAP3 S_PMAP5 S_PMAP6 THUSTR_12 "level 12: crater" HUSTR_7 "level 7: dead simple" ST_POSITIVE weapontype_t viewactive divline_t key_map_east key_prevweapon STSTR_MUS "Music Change" GOTHTHBONUS "Picked up a health bonus." VIEWHEIGHT (41*FRACUNIT) SPR_BFE1 SPR_BFE2 ds_source maxx KEY_UPARROW 0xad pendingweapon PHUSTR_13 "level 13: the crypt" S_RTORCHSHRT2 S_RTORCHSHRT3 S_RTORCHSHRT4 S_CHAINUP SPR_BFUG S_TROO_PAIN downstate AMSTR_MARKSCLEARED "All Marks Cleared" nexttic specialdata SPR_BON1 SPR_BON2 key_usehealth PHUSTR_21 "level 21: slayer" PT_ADDTHINGS 2 S_SKEL_DIE2 doom1_endmsg S_PLAY_DIE7 bprev AM_updateLightLev S_YKEY S_SSWV_PAIN2 HUSTR_KEYGREEN 'g' va_start(v,l) __builtin_va_start(v,l) HUSTR_E4M6 "E4M6: Against Thee Wickedly" S_HEARTCOL GREENRANGE 16 NET_MAXPLAYERS 8 S_SSWV_ATK1 S_SSWV_ATK2 S_SSWV_ATK3 S_SSWV_ATK4 S_SSWV_ATK5 S_SSWV_ATK6 screenheightarray S_TECH2LAMP4 S_SOUL SPR_BFGF SPR_BFGG S_SPOS_DIE1 S_SPOS_DIE2 S_SPOS_DIE3 S_SPOS_DIE4 S_SPOS_DIE5 __D_THINK__  SPR_TFOG tmfloorz MSGON "Messages ON" spritetopoffset S_SKULL_DIE1 S_SKULL_DIE2 S_SKULL_DIE3 S_SKULL_DIE4 SCREENHEIGHT_4_3 240 key_weapon2 key_weapon3 key_weapon4 key_weapon5 key_weapon6 key_weapon7 key_weapon8 DEH_STR_H  S_SKEL_RUN1 S_SKEL_RUN2 S_SKEL_RUN3 S_SKEL_RUN4 S_SKEL_RUN5 S_SKEL_RUN6 S_SKEL_RUN7 S_SKEL_RUN8 S_SKEL_RUN9 S_SMOKE3 C2TEXT "YOU HAVE WON! YOUR VICTORY HAS ENABLED\n" "HUMANKIND TO EVACUATE EARTH AND ESCAPE\n""THE NIGHTMARE.  NOW YOU ARE THE ONLY\n""HUMAN LEFT ON THE FACE OF THE PLANET.\n""CANNIBAL MUTATIONS, CARNIVOROUS ALIENS,\n""AND EVIL SPIRITS ARE YOUR ONLY NEIGHBORS.\n""YOU SIT BACK AND WAIT FOR DEATH, CONTENT\n""THAT YOU HAVE SAVED YOUR SPECIES.\n""\n""BUT THEN, EARTH CONTROL BEAMS DOWN A\n""MESSAGE FROM SPACE: \"SENSORS HAVE LOCATED\n""THE SOURCE OF THE ALIEN INVASION. IF YOU\n""GO THERE, YOU MAY BE ABLE TO BLOCK THEIR\n""ENTRY.  THE ALIEN BASE IS IN THE HEART OF\n""YOUR OWN HOME CITY, NOT FAR FROM THE\n""STARPORT.\" SLOWLY AND PAINFULLY YOU GET\n""UP AND RETURN TO THE FRAY." KEY_STRAFE_L 0xa0 raiseToNearestAndChange GOTCLIPBOX "Picked up a box of bullets." S_CPOS_RAISE4 S_HEAD_DIE1 S_HEAD_DIE2 S_HEAD_DIE3 S_HEAD_DIE5 S_HEAD_DIE6 SPR_SMBT S_SKULL_RUN2 menuactive GOTARMOR "Picked up the armor." thinkercap SLOPEBITS 11 NUMCARDS MTF_AMBUSH 8 key_map_zoomin key_lookdown S_BSPI_DIE2 THINGCOLORS GREENS S_BSPI_DIE3 KEY_RIGHTARROW 0xae S_BSPI_DIE4 S_BSPI_DIE5 S_PLAY_PAIN S_BSPI_DIE6 S_PISTOLFLASH key_arti_blastradius S_DEADSTICK it_redskull SPR_CLIP __R_MAIN__  STSTR_CLEV "Changing Level..." S_DSGUN1 ANG60 (ANG180 / 3) key_arti_teleportother exe_hacx LOADNET "you can't do load while in a net game!\n\n"PRESSKEY cheating intercept_t numnodes MT_KEEN S_PSTR S_COMMKEEN2 S_COMMKEEN3 S_COMMKEEN4 S_COMMKEEN5 S_COMMKEEN6 S_COMMKEEN7 S_COMMKEEN8 ST_WIDTH SCREENWIDTH S_SPAWNFIRE2 SPR_BOSF AM_NUMMARKPOINTS 10 SPR_BOSS S_SHEL AM_clearMarks SPR_POL1 SPR_POL2 SPR_POL5 SPR_POL6 SPR_FSKU KEY_F12 (0x80+0x58) uint8_t SPR_CAND statenum_t S_CPOS_XDIE1 S_CPOS_XDIE2 S_CPOS_XDIE3 S_PLAS S_CPOS_XDIE5 S_CPOS_XDIE6 S_KEENSTND S_PLAY mpoint_t CXMTOF(x) (f_x + MTOF((x)-m_x)) PRESSYN "press y or n." S_FATT_DIE7 S_FATT_DIE8 THUSTR_22 "level 22: habitat" PHUSTR_20 "level 20: the death domain" __R_BSP__  KEY_TAB 9 S_GTORCHSHRT sprtopscreen S_BOS2_STND SPR_SARG PD_YELLOWO "You need a yellow key to activate this object" pack_tnt am_clip HUSTR_CHATMACRO0 "No" USERANGE (64*FRACUNIT) sidedef S_BLOOD1 opentop startepisode S_BKEY S_POSS_STND mceilingclip KEY_LEFTARROW 0xac M_ZOOMIN ((int) (1.02*FRACUNIT)) __R_SEGS__  dc_colormap precache viewx viewy viewz float S_CYBER_RUN1 S_CYBER_RUN3 S_CYBER_RUN4 S_CYBER_RUN5 S_CYBER_RUN6 S_CYBER_RUN7 S_CYBER_RUN8 param_chars_read SPR_SMGT PLATWAIT 3 SPR_PINS S_FLOATSKULL2 S_FLOATSKULL3 HUSTR_TALKTOSELF2 "Who's there?" PHUSTR_28 "level 28: the sewers" SPR_VILE S_BFGEXP AM_LevelInit mouse_acceleration S_BTORCHSHRT4 HUSTR_9 "level 9: the pit" P2TEXT "Even the deadly Arch-Vile labyrinth could\n""not stop you, and you've gotten to the\n""prototype Accelerator which is soon\n""efficiently and permanently deactivated.\n""\n""You're good at that kind of thing." CC_PAIN "PAIN ELEMENTAL" HUSTR_MSGU "[Message unsent]" PHUSTR_16 "level 16: the omen" S_BOS2_STND2 S_SGUN1 S_SGUN2 S_SGUN3 S_SGUN4 S_SGUN5 S_SGUN6 S_SGUN7 S_SGUN8 S_SGUN9 FDWALLRANGE BROWNRANGE SECRETWALLCOLORS WALLCOLORS S_MEDI S_SARG_PAIN2 tantoangle S_VILE_STND DETAILHI "High detail" SPR_TGRN ev_joystick rw_stopx cheat_mypos lightlevel f_oldloc MT_HEADSHOT wbplayerstruct_t floatok SPR_SMIT S_BSPI_RAISE4 S_SKULLCOL SPR_SKUL startloadgame key_menu_down usedown sk_baby S_SSWV_DIE1 S_SSWV_DIE2 S_SSWV_DIE3 S_SSWV_DIE4 S_SSWV_DIE5 SPR_TROO KEYP_0 0 S_BOS2_ATK1 S_BOS2_ATK2 S_BOS2_ATK3 S_SKEL_RAISE1 S_SKEL_RAISE2 S_SKEL_RAISE3 S_SKEL_RAISE4 S_SKEL_RAISE5 S_SKEL_RAISE6 PHUSTR_8 "level 8: realm" mousebstraferight S_BAR2 MT_EXTRABFG degenmobj_t SPR_AMMO pw_invisibility BLACK 0 GOTBLUECARD "Picked up a blue keycard." S_CANDELABRA S_POSS_ATK1 S_POSS_ATK2 S_POSS_ATK3 PHUSTR_26 "level 26: bunker" PHUSTR_5 "level 5: ghost town" S_TROO_XDIE1 S_TROO_XDIE2 S_TROO_XDIE3 S_TROO_XDIE4 key_invquery ev_keyup S_TROO_XDIE8 HUSTR_18 "level 18: the courtyard" KEY_HOME (0x80+0x47) __R_LOCAL__  MT_SMOKE st_backing_screen MLIBC_POSIX_STRING_H  key_menu_activate S_MEGA KEY_F5 (0x80+0x3f) GS_DEMOSCREEN SPR_CYBR ANG270 0xc0000000 THUSTR_9 "level 9: stronghold" SPR_SBOX SPR_POSS SPR_BFS1 key_menu_screenshot SPR_IFOG S_BLOODYTWITCH3 S_BLOODYTWITCH4 PD_BLUEK "You need a blue key to open this door" YELLOWRANGE 1 wad_file_class_t subsector joybstraferight S_SSWV_XDIE2 KEY_USE 0xa2 FEATURE_SOUND texturetranslation PD_YELLOWK "You need a yellow key to open this door" drawseg_t THUSTR_13 "level 13: nukage processing" GOTCELLBOX "Picked up an energy cell pack." P3TEXT "You've bashed and battered your way into\n""the heart of the devil-hive.  Time for a\n""Search-and-Destroy mission, aimed at the\n""Gatekeeper, whose foul offspring is\n""cascading to Earth.  Yeah, he's bad. But\n""you know who's worse!\n""\n""Grinning evilly, you check your gear, and\n""get ready to give the bastard a little Hell\n""of your own making!" maxsecret wp_missile S_VILE_ATK1 S_VILE_ATK2 S_VILE_ATK3 S_VILE_ATK4 nextstate S_VILE_ATK6 S_VILE_ATK7 S_VILE_ATK8 S_VILE_ATK9 GAMMALVL1 "Gamma correction level 1" S_SPOS_STND2 va_arg(v,l) __builtin_va_arg(v,l) S_RKEY2 S_SPID_PAIN STSTR_BEHOLD "inVuln, Str, Inviso, Rad, Allmap, or Lite-amp" THUSTR_19 "level 19: shipping/respawning" HUSTR_KEYRED 'r' ceilingpic S_SSWV_PAIN am_shell SIL_BOTH 3 MAXLIGHTZ 128 PHUSTR_22 "level 22: impossible mission" mobjinfo_t firstflat NUMSTATES seestate mtof_zoommul S_SHOT S_COMMKEEN9 LIGHTZSHIFT 20 fpoint_t MT_CHAINGUY HUSTR_E1M7 "E1M7: Computer Station" MT_KNIGHT S_BFGUP ticdup S_HEAD_PAIN2 S_HEAD_PAIN3 CC_HEAVY "HEAVY WEAPON DUDE" key_map_follow S_SARG_RAISE1 S_SARG_RAISE2 S_SARG_RAISE3 S_SARG_RAISE4 S_SARG_RAISE5 S_SARG_RAISE6 E4TEXT "the spider mastermind must have sent forth\n""its legions of hellspawn before your\n""final confrontation with that terrible\n""beast from hell.  but you stepped forward\n""and brought forth eternal damnation and\n""suffering upon the horde as a true hero\n""would in the face of something so evil.\n""\n""besides, someone was gonna pay for what\n""happened to daisy, your pet rabbit.\n""\n""but now, you see spread before you more\n""potential pain and gibbitude as a nation\n""of demons run amok among our cities.\n""\n""next stop, hell on earth!" GameVersion_t S_RSKULL2 S_BOSS_PAIN2 THINGRANGE GREENRANGE ammotype_t key_lookup musicVolume S_SSWV_RUN4 S_BON1A S_BON1B MT_TFOG S_BON1D S_BON1E joybjump viewangletox attacksound SAVEDEAD "you can't save if you aren't playing!\n\n"PRESSKEY respawnmonsters ENDGAME "are you sure you want to end the game?\n\n"PRESSYN gamemode FLOATSPEED (FRACUNIT*4) key_map_toggle S_ROCK S_BON2C S_BON2D S_BON2E angle_t KEY_PGDN (0x80+0x51) gamemission spriteoffset weaponinfo_t viewsin S_TECHLAMP3 S_DSGUNFLASH1 S_HANGTNOBRAIN S_PAIN_PAIN2 M_snprintf S_PUNCHDOWN file_class S_TRACEEXP2 KEYP_EQUALS KEY_EQUALS S_HEAD_RAISE1 S_HEAD_RAISE2 S_HEAD_RAISE3 S_HEAD_RAISE4 lastlevel key_multi_msg PHUSTR_15 "level 15: the twilight" PU_CACHE max_x max_y MAPBLOCKSIZE (MAPBLOCKUNITS*FRACUNIT) __D_LOOP__  __M_CHEAT__  SPR_COL2 leveljuststarted meleestate __DOOMDEF__  S_MISSILEFLASH2 S_MISSILEFLASH4 S_CYBER_STND2 MT_CLIP __R_DATA__  PHUSTR_19 "level 19: nme" S_SKULL_RUN1 indetermined perpetualRaise S_LIGHTDONE _VA_LIST_  HUSTR_19 "level 19: the citadel" wp_nochange S_SPID_RUN10 S_SPID_RUN11 S_SPID_RUN12 S_SARG_PAIN THUSTR_3 "level 3: power control" MT_BOSSTARGET MT_TELEPORTMAN NET_TICDIFF_TURN (1 << 2) S_TFOG2 S_TFOG3 S_TFOG4 S_TFOG5 S_TFOG6 S_TFOG7 S_TFOG8 S_TFOG9 S_POSS_PAIN2 markceiling S_SPAWNFIRE8 curline S_BOS2_DIE1 S_BOS2_DIE2 S_BOS2_DIE3 S_BOS2_DIE4 S_BOS2_DIE5 S_BOS2_DIE6 S_BOS2_DIE7 SPR_BSKU singletics BUTTONTIME 35 HUSTR_CHATMACRO7 "Come here!" silentCrushAndRaise S_REDTORCH2 S_REDTORCH3 S_REDTORCH4 S_TALLGRNCOL S_BFGFLASH1 S_BFGFLASH2 S_REDTORCH S_POSS_DIE1 S_POSS_DIE2 S_POSS_DIE3 S_PISTOLUP S_POSS_DIE5 key_menu_incscreen S_PLASEXP5 S_BPAK ML_SOUNDBLOCK 64 GRIDCOLORS (GRAYS + GRAYSRANGE/2) spritewidth MAXSPECIALCROSS 20 pspriteiscale S_VILE_ATK10 spritenum_t snd_SfxDevice HUSTR_15 "level 15: industrial zone" HUSTR_23 "level 23: barrels o' fun" cheat_mus FASTDARK 15 S_EXPLODE1 S_EXPLODE2 S_EXPLODE3 netcmds __R_DEFS__  MAX_MOUSE_BUTTONS 8 ds_p SPR_HDB1 SPR_HDB2 SPR_HDB3 SPR_HDB4 SPR_HDB5 SPR_HDB6 ds_y plyr S_FIRE3 S_BOSS_RUN1 S_BOSS_RUN2 S_BOSS_RUN3 S_BOSS_RUN4 S_BOSS_RUN5 S_BOSS_RUN6 S_BOSS_RUN7 S_BOSS_RUN8 misc1 misc2 __SHA1_H__  KEY_F10 (0x80+0x44) ST_NEGATIVE P1TEXT "You gloat over the steaming carcass of the\n""Guardian.  With its death, you've wrested\n""the Accelerator from the stinking claws\n""of Hell.  You relax and glance around the\n""room.  Damn!  There was supposed to be at\n""least one working prototype, but you can't\n""see it. The demons must have taken it.\n""\n""You must find the prototype, or all your\n""struggles will have been wasted. Keep\n""moving, keep fighting, keep killing.\n""Oh yes, keep living, too." st_notify S_BRBALLX1 S_BRBALLX2 markfloor S_SKEL_STND HUSTR_12 "level 12: the factory" PD_REDO "You need a red key to activate this object" linedef basedefault KEY_F6 (0x80+0x40) S_FATT_RUN1 S_FATT_RUN2 S_FATT_RUN4 S_FATT_RUN5 S_FATT_RUN6 MT_VILE S_FATT_DIE6 S_FATT_RUN9 SPR_FCAN mousebfire key_map_south S_VILE_DIE3 S_VILE_DIE4 S_VILE_DIE5 S_VILE_DIE6 S_BRAINEXPLODE1 S_BRAINEXPLODE2 S_BRAINEXPLODE3 S_CHAINDOWN S_YKEY2 KEY_NUMLOCK (0x80+0x45) HUSTR_16 "level 16: suburbs" CC_CACO "CACODEMON" AM_MSGHEADER (('a'<<24)+('m'<<16)) vscalelight ds_x1 ds_x2 PHUSTR_6 "level 6: baron's lair" wbstartstruct_t AM_saveScaleAndLoc S_TRACEEXP1 CHEAT(value,parameters) { value, sizeof(value) - 1, parameters, 0, 0, "" } S_TRACEEXP3 KEYP_9 KEY_PGUP fixed_t S_SUIT HUSTR_CHATMACRO5 "You suck!" mouse_threshold key_menu_save snext S_VILE_DIE10 maxfrags byte fuzzcolfunc S_CELL HUSTR_E4M7 "E4M7: And Hell Followed" NET_TICDIFF_STRIFE (1 << 7) GOTARMBONUS "Picked up an armor bonus." S_CPOS_RUN1 S_CPOS_RUN2 S_CPOS_RUN3 S_CPOS_RUN4 S_CPOS_RUN5 S_CPOS_RUN6 S_CPOS_RUN7 S_CPOS_RUN8 GRAVITY FRACUNIT joybuse SPR_BSPI S_TFOG01 S_TFOG02 S_SPAWN4 DOOM_VERSION 109 cheat_clev SPR_SMRT PHUSTR_24 "level 24: the final frontier" ceilingheight MAXMOVE (30*FRACUNIT) activeceilings V_DrawPatch S_CANDLESTIK AM_doFollowPlayer crushAndRaise HUSTR_KEYINDIGO 'i' key_menu_left S_SKULL_STND2 QSPROMPT "quicksave over your game named\n\n'%s'?\n\n"PRESSYN rw_distance S_TFOG10 PD_REDK "You need a red key to open this door" HUSTR_CHATMACRO9 "Yes" ps_weapon DOOM_FEATURES_H  sk_nightmare S_RTORCHSHRT SPR_CELL SPR_CELP LINE_NEVERSEE ML_DONTDRAW S_BFGSHOT _VA_LIST_T_H  statusbaractive KEY_RALT (0x80+0x38) devparm key_map_grid m_x2 MT_SKULL pack_chex GOTCHAINGUN "You got the chaingun!" S_PINV4 last numsectors SPR_MANF S_BLUETORCH gammatable S_SARG_RUN3 _wad_file_s HUSTR_E3M9 "E3M9: Warrens" HUSTR_PLRRED "Red: " SPR_SMT2 SPR_RKEY THUSTR_17 "level 17: processing area" marknums painstate S_CYBER_STND HUSTR_E1M3 "E1M3: Toxin Refinery" HUSTR_E2M8 "E2M8: Tower of Babel" numsegs AM_drawThings mline_t KEYP_MULTIPLY '*' S_SPOS_RUN6 am_cell movedir HUSTR_8 "level 8: tricks and traps" S_SPOS_RUN8 THUSTR_4 "level 4: wormhole" S_FATT_DIE10 MT_IFOG missilestate max_h exe_doom_1_666 KEY_PGUP (0x80+0x49) tmceilingz SPR_HEAD MT_PLASMA HUSTR_32 "level 32: grosse" C5TEXT "CONGRATULATIONS, YOU'VE FOUND THE SECRET\n""LEVEL! LOOKS LIKE IT'S BEEN BUILT BY\n""HUMANS, RATHER THAN DEMONS. YOU WONDER\n""WHO THE INMATES OF THIS CORNER OF HELL\n""WILL BE." SIL_TOP 2 SPR_FATB SECRETWALLRANGE WALLRANGE SPR_FATT YELLOWS (256-32+7) __DOOMDATA__  S_TECHLAMP KEYP_PERIOD 0 pw_strength PHUSTR_23 "level 23: tombstone" soundtarget gameepisode mousebuse respawnparm CEILSPEED FRACUNIT outside __I_TIMER__  HUSTR_26 "level 26: the abandoned mines" S_HANGTLOOKDN key_pause BLUERANGE 8 backpack S_ARACH_PLAZ2 SPR_YKEY MT_SPIDER gameskill S_SMALLPOOL options sprnames GGSAVED "game saved." THUSTR_16 "level 16: deepest reaches" CC_MANCU "MANCUBUS" iquetail S_CYBER_ATK1 S_CYBER_ATK2 S_CYBER_ATK3 S_CYBER_ATK4 S_CYBER_ATK5 S_CYBER_ATK6 KEY_PAUSE 0xff S_VILE_DIE1 doom2_endmsg THUSTR_24 "level 24: quarry" S_BIGTREE SPR_SOUL ds_xstep SPR_CPOS NEWGAME "you can't start a new game\n""while in a network game.\n\n"PRESSKEY numsides distscale S_PINV2 S_PINV3 MT_FATSO HUSTR_CHATMACRO2 "I'm OK." button_t S_SSWV_STND2 PHUSTR_10 "level 10: onslaught" outcode2 S_POSS_XDIE4 SPR_PUFF S_POSS_XDIE6 S_POSS_XDIE8 SPR_TLMP S_FLOATSKULL AM_MSGENTERED (AM_MSGHEADER | ('e'<<8)) key_map_west ANG_MAX 0xffffffff DETAILLO "Low detail" S_SPOS_PAIN cheat_amap REDS (256-5*16) S_BFGSHOT2 NET_TICDIFF_BUTTONS (1 << 3) S_SKULL_PAIN key_down DOOM_191_VERSION 111 S_HANGNOGUTS vanilla_keyboard_mapping litelevels linetarget key_demo_quit MAXVISSPRITES 128 STSTR_DQDON "Degreelessness Mode On" cheat_commercial_noclip numvertexes PST_REBORN shareware PU_NUM_TAGS S_COMMKEEN min_x none S_BAR1 MAXPLAYERNAME 30 rw_x S_HEAD_PAIN MT_CYBORG PU_PURGELEVEL spriteframes spritedef_t S_SKEL_DIE1 S_SKEL_DIE3 S_SKEL_DIE4 SPR_PSTR S_SKEL_DIE6 MAXNETNODES 16 hexen P6TEXT "Betcha wondered just what WAS the hardest\n""level we had ready for ya?  Now you know.\n""No one gets out alive." MT_MISC31 S_LAUN SPR_TLP2 key_arti_health MT_MISC37 wp_chainsaw SPR_BAL1 SPR_BAL2 SPR_SHEL snd_DesiredMusicDevice SPR_BAL7 V_PATCH_H  BASETHRESHOLD 100 PHUSTR_12 "level 12: speed" CC_CYBER "THE CYBERDEMON" GOTCLIP "Picked up a clip." btimer screen_width itemrespawnque S_TROO_RAISE1 S_TROO_RAISE2 S_TROO_RAISE3 S_TROO_RAISE4 S_TROO_RAISE5 S_MGUN SPR_PLAY ANG180 0x80000000 backsector MTF_HARD 4 lowerAndCrush GOTREDCARD "Picked up a red keycard." silhouette S_BFGLAND plattype_e MT_CHAINGUN KEYP_1 KEY_END T6TEXT "Time for a vacation. You've burst the\n""bowels of hell and by golly you're ready\n""for a break. You mutter to yourself,\n""Maybe someone else can kick Hell's ass\n""next time around. Ahead lies a quiet town,\n""with peaceful flowing water, quaint\n""buildings, and presumably no Hellspawn.\n""\n""As you step off the transport, you hear\n""the stomp of a cyberdemon's iron shoe." MT_ROCKET GOTLAUNCHER "You got the rocket launcher!" S_HEARTCOL2 MT_MISC44 MT_MISC45 HUSTR_E4M9 "E4M9: Fear" MT_MISC47 validcount S_VILE_HEAL3 ML_SECRET 32 THUSTR_32 "level 32: caribbean" FTOM(x) FixedMul(((x)<<16),scale_ftom) deathmatch_p HUSTR_4 "level 4: the focus" KEYP_3 KEY_PGDN SPR_CEYE THUSTR_28 "level 28: heck" E3TEXT "The loathsome spiderdemon that\n""masterminded the invasion of the moon\n""bases and caused so much death has had\n""its ass kicked for all time.\n""\n""A hidden doorway opens and you enter.\n""You've proven too tough for Hell to\n""contain, and now Hell at last plays\n""fair -- for you emerge from the door\n""to see the green fields of Earth!\n""Home at last.\n" "\n""You wonder what's been happening on\n""Earth while you were battling evil\n""unleashed. It's good that no Hell-\n""spawn could have come through that\n""door with you ..." F_PANINC 4 S_CHAIN STSTR_CHOPPERS "... doesn't suck - GM" bsilheight KEY_ENTER 13 children textureoffset MAX_CHEAT_LEN 25 AM_MSGEXITED (AM_MSGHEADER | ('x'<<8)) AM_getIslope S_TECH2LAMP2 S_TECH2LAMP3 S_PAIN_RUN1 S_PAIN_RUN2 S_PAIN_RUN3 S_PAIN_RUN4 S_PAIN_RUN5 S_PAIN_RUN6 S_FATT_DIE3 S_FATT_DIE4 S_SMOKE1 S_SMOKE2 S_BEXP S_SMOKE4 S_SMOKE5 S_PISTOL2 skyflatnum S_FATT_DIE9 MAXPLAYERS 4 totalsecret ceilingplane MT_MISC51 S_DSNR2 cheat_ammonokey S_SPOS_PAIN2 S_PUNCHUP RANGECHECK  S_SKEL_RUN10 S_SKEL_RUN11 S_SKEL_RUN12 reactiontime SPR_MEDI maxitems S_BFGDOWN openbottom NET_TICDIFF_CONSISTANCY (1 << 4) __R_DRAW__  S_BRBALLX3 spriteframe_t thintriangle_guy ML_MAPPED 256 S_BSPI_RAISE6 S_BRAIN_DIE2 S_BRAIN_DIE3 S_BRAIN_DIE4 crush STSTR_NCOFF "No Clipping Mode OFF" ANGLETOFINESHIFT 19 SPR_PAIN wminfo S_SAW1 S_SAW2 S_SAW3 S_HEADCANDLES2 bmapheight MT_SUPERSHOTGUN C1TEXT "YOU HAVE ENTERED DEEPLY INTO THE INFESTED\n" "STARPORT. BUT SOMETHING IS WRONG. THE\n" "MONSTERS HAVE BROUGHT THEIR OWN REALITY\n" "WITH THEM, AND THE STARPORT'S TECHNOLOGY\n" "IS BEING SUBVERTED BY THEIR PRESENCE.\n" "\n""AHEAD, YOU SEE AN OUTPOST OF HELL, A\n" "FORTIFIED ZONE. IF YOU CAN GET PAST IT,\n" "YOU CAN PENETRATE INTO THE HAUNTED HEART\n" "OF THE STARBASE AND FIND THE CONTROLLING\n" "SWITCH WHICH HOLDS EARTH'S POPULATION\n" "HOSTAGE." xdeathstate S_CYBER_DIE1 S_CYBER_DIE2 S_CYBER_DIE3 S_CYBER_DIE4 S_CYBER_DIE5 S_CYBER_DIE6 S_CYBER_DIE7 S_CYBER_DIE8 S_CYBER_DIE9 SWSTRING "this is the shareware version of doom.\n\n""you need to order the entire trilogy.\n\n"PRESSKEY MT_FATSHOT MT_BABY V_MarkRect mobjflags picnum SPR_BAR1 retail S_TRACER S_GREENTORCH position didsecret S_HEAD_RAISE5 old_m_x MT_SPAWNSHOT S_SPID_RUN1 S_SPID_RUN2 S_FATT_STND S_BRAIN S_SPID_ATK1 S_SPID_RUN6 S_FIRE10 S_FIRE11 S_FIRE12 S_FIRE13 S_FIRE14 S_FIRE15 S_FIRE16 S_FIRE17 S_FIRE18 S_FIRE19 S_BSPI_DIE7 BROWNRANGE 16 SPR_MEGA HUSTR_CHATMACRO1 "I'm ready to kick butt!" GRIDRANGE 0 bodyqueslot activesound wp_shotgun killcount HUSTR_20 "level 20: gotcha!" MT_MISC71 HUSTR_21 "level 21: nirvana" followplayer HUSTR_30 "level 30: icon of sin" S_ARACH_PLEX3 ceilingfunc_t S_FIRE20 S_FIRE21 S_FIRE22 S_FIRE23 S_FIRE24 S_FIRE25 S_FIRE26 S_FIRE27 S_FIRE28 S_FIRE29 PRESSKEY "press a key." S_DSGUN2 S_DSGUN3 S_DSGUN4 S_DSGUN5 S_DSGUN6 S_DSGUN7 S_DSGUN8 S_DSGUN9 DEH_VANILLA_NUMSTATES 966 CC_ARACH "ARACHNOTRON" LIGHTLEVELS 16 __DSTRINGS__  NUMCOLORMAPS 32 ONFLOORZ INT_MIN sk_easy ceilingline STSTR_DQDOFF "Degreelessness Mode Off" their_colors NF_SUBSECTOR 0x8000 S_FIRE30 ev_mouse PHUSTR_29 "level 29: odyssey of noises" namebuf GRAYS (6*16) S_TRACER2 QUITMSG "are you sure you want to\nquit this great game?" projection ANG90 0x40000000 S_SPAWN1 S_SPAWN2 S_SPAWN3 cheat_ammo S_BROK S_SSWV_RAISE1 MT_MISC80 S_PUFF1 S_PUFF3 S_PUFF4 __va_list__  acp1 acp2 PST_DEAD YOURCOLORS WHITE PHUSTR_32 "level 32: go 2 it" SPR_SHOT FEATURE_MULTIPLAYER pw_infrared screensaver_mode GAMMALVL4 "Gamma correction level 4" HUSTR_E2M9 "E2M9: Fortress of Mystery" S_BOSS_ATK1 S_BOSS_ATK2 S_BOSS_ATK3 key_menu_detail mfloorclip mousebstrafe S_SAWDOWN tracer key_fire buttonlist GOTMEDIKIT "Picked up a medikit." startskill GOTVISOR "Light Amplification Visor" S_FATT_ATK1 S_FATT_ATK2 S_FATT_ATK3 S_FATT_ATK4 S_FATT_ATK5 S_FATT_ATK6 S_FATT_ATK7 S_FATT_ATK8 S_FATT_ATK9 mobjinfo S_HANGTLOOKUP HUSTR_E3M4 "E3M4: House of Pain" GOTSHELLBOX "Picked up a box of shotgun shells." AM_drawCrosshair S_PLASEXP HUSTR_E3M5 "E3M5: Unholy Cathedral" S_SKULL_ATK2 GOTSHOTGUN2 "You got the super shotgun!" HUSTR_13 "level 13: downtown" slopetype_t MT_PUFF PHUSTR_1 "level 1: congo" T4TEXT "Suddenly, all is silent, from one horizon\n""to the other. The agonizing echo of Hell\n""fades away, the nightmare sky turns to\n""blue, the heaps of monster corpses start \n""to evaporate along with the evil stench \n""that filled the air. Jeeze, maybe you've\n""done it. Have you really won?\n""\n""Something rumbles in the distance.\n""A blue light begins to glow inside the\n""ruined skull of the demon-spitter." SPR_ROCK parameter_buf GOTCELL "Picked up an energy cell." isaline olddirection S_BSPI_RUN2 S_BSPI_RUN3 S_BSPI_RUN4 S_BSPI_RUN5 S_BSPI_RUN6 S_BSPI_RUN7 S_BSPI_RUN8 S_BSPI_RUN9 SPR_BLUD lowres_turn MT_BRUISERSHOT MISSILERANGE (32*64*FRACUNIT) dc_x spawnhealth CEILWAIT 150 GS_FINALE S_CPOS_ATK1 S_CPOS_ATK2 S_CPOS_ATK3 S_CPOS_ATK4 forwardmove key_map_zoomout fixedcolormap S_BLOODYTWITCH cheatseq_t rejectmatrix min_h epsd SPR_FIRE firstspritelump loopcount S_PINS3 timelimit aspect_ratio_correct key_left S_TALLREDCOL linecount itemrespawntime SPR_PINV PU_STATIC S_CPOS_STND HUSTR_E3M1 "E3M1: Hell Keep" S_SKEL_FIST2 __D_ITEMS__  modifiedgame MT_MISC0 MT_MISC1 MT_MISC2 MT_MISC3 MT_MISC4 MT_MISC5 MT_MISC6 S_SKULL_ATK1 S_BRBALL1 S_BRBALL2 S_SKULL_ATK3 scaledviewwidth detailshift GOTYELWSKUL "Picked up a yellow skull key." CC_IMP "IMP" viewcos SPR_SHT2 PLAYERRADIUS 16*FRACUNIT ds_ystep THUSTR_11 "level 11: storage facility" SPR_SHTF SPR_SHTG S_BON2 PHUSTR_9 "level 9: abattoire" MT_UNDEAD S_TROO_RUN1 S_TROO_RUN2 S_TROO_RUN3 S_TROO_RUN4 S_TROO_RUN5 S_TROO_RUN6 S_TROO_RUN7 S_TROO_RUN8 _ANSI_STDARG_H_  S_BSPI_RUN1 pad2 pad3 DOOUTCODE(oc,mx,my) (oc) = 0; if ((my) < 0) (oc) |= TOP; else if ((my) >= f_h) (oc) |= BOTTOM; if ((mx) < 0) (oc) |= LEFT; else if ((mx) >= f_w) (oc) |= RIGHT; lineguylines __D_ENGLSH__  INITSCALEMTOF (.2*FRACUNIT) S_COLU SPR_ELEC S_VILE_RUN1 dclick_use S_VILE_RUN2 S_KEENPAIN ML_BLOCKMONSTERS 2 HUSTR_PLRBROWN "Brown: " DBITS (FRACBITS-SLOPEBITS) S_SKULL_PAIN2 seesound S_CYBER_RUN2 AM_drawFline AMSTR_GRIDON "Grid ON" SPR_BPAK XHAIRCOLORS GRAYS S_ARACH_PLEX2 key_speed S_ARACH_PLEX4 S_ARACH_PLEX5 S_COMMKEEN10 S_BOS2_PAIN lighttable_t CENTERY (SCREENHEIGHT/2) HUSTR_31 "level 31: wolfenstein" NETEND "you can't end a netgame!\n\n"PRESSKEY max_w vissprite_p S_SPID_DIE10 S_SPID_DIE11 S_POSS_PAIN AM_activateNewScale GOTMSPHERE "MegaSphere!" DOSY "(press y to quit to dos.)" S_GREENTORCH2 S_GREENTORCH3 S_GREENTORCH4 KEYP_ENTER KEY_ENTER MTF_NORMAL 2 cheat_god GOTBFG9000 "You got the BFG9000!  Oh, yes." DEH_AddStringReplacement(x,y)  where C4TEXT "THE HORRENDOUS VISAGE OF THE BIGGEST\n""DEMON YOU'VE EVER SEEN CRUMBLES BEFORE\n""YOU, AFTER YOU PUMP YOUR ROCKETS INTO\n""HIS EXPOSED BRAIN. THE MONSTER SHRIVELS\n""UP AND DIES, ITS THRASHING LIMBS\n""DEVASTATING UNTOLD MILES OF HELL'S\n""SURFACE.\n""\n""YOU'VE DONE IT. THE INVASION IS OVER.\n""EARTH IS SAVED. HELL IS A WRECK. YOU\n""WONDER WHERE BAD FOLKS WILL GO WHEN THEY\n""DIE, NOW. WIPING THE SWEAT FROM YOUR\n""FOREHEAD YOU BEGIN THE LONG TREK BACK\n""HOME. REBUILDING EARTH OUGHT TO BE A\n""LOT MORE FUN THAN RUINING IT WAS.\n" S_PISTOL1 S_PISTOL3 S_PISTOL4 exe_strife_1_31 SPR_PLSE SPR_PLSF SPR_PLSG cheat_powerup FEATURE_DEHACKED SPR_PLSS DEH_fprintf fprintf DEH_snprintf snprintf HUSTR_27 "level 27: monster condo" diskicon_readbytes blockmap GLOWSPEED 8 S_SSWV_XDIE1 S_SSWV_XDIE3 S_SSWV_XDIE4 S_PAIN_RAISE1 S_PAIN_RAISE2 S_PAIN_RAISE3 S_PAIN_RAISE4 S_PAIN_RAISE5 S_PAIN_RAISE6 S_DEADBOTTOM CDWALLCOLORS YELLOWS SPR_SUIT ps_flash key_arti_poisonbag autostart __D_MODE__  S_PLAY_RUN1 S_PLAY_RUN2 S_PLAY_RUN3 S_PLAY_RUN4 S_BOSS_STND2 ANG45 0x20000000 numsubsectors S_VILE_PAIN key_menu_abort S_IFOG2 S_IFOG3 S_IFOG4 S_IFOG5 bonuscount S_BOSS_DIE1 S_BOSS_DIE2 S_BOSS_DIE3 S_BOSS_DIE5 S_BOSS_DIE6 S_BOSS_DIE7 MT_PLAYER S_HEADONASTICK finesine S_CPOS_XDIE4 key_invkey segtextured AM_findMinMaxBoundaries S_SSWV_RAISE2 S_SSWV_RAISE3 S_SSWV_RAISE4 S_SSWV_RAISE5 HUSTR_E2M5 "E2M5: Command Center" S_POSS_XDIE1 S_POSS_XDIE2 S_POSS_XDIE3 S_POSS_XDIE5 show_diskicon S_POSS_XDIE7 DEH_printf printf S_POSS_XDIE9 ML_DONTDRAW 128 BACKGROUND BLACK S_SPOS_RUN3 S_SPOS_RUN5 cheat_noclip joybstrafeleft GameMission_t visplane_t SPR_SSWV P4TEXT "The Gatekeeper's evil face is splattered\n""all over the place.  As its tattered corpse\n""collapses, an inverted Gate forms and\n""sucks down the shards of the last\n""prototype Accelerator, not to mention the\n""few remaining demons.  You're done. Hell\n""has gone back to pounding bad dead folks \n""instead of good live ones.  Remember to\n""tell your grandkids to put a rocket\n""launcher in your coffin. If you go to Hell\n""when you die, you'll need it for some\n""final cleaning-up ..." S_PLASEXP2 S_PLASEXP3 S_PLASEXP4 S_CHAIN1 S_CHAIN2 S_CHAIN3 S_PLAY_PAIN2 sk_medium S_FIRE8 centeryfrac MT_MEGA bmapwidth NUMPSPRITES joybprevweapon tinttable usegamma dscalelight HUSTR_14 "level 14: the inmost dens" S_EVILEYE2 S_EVILEYE3 S_EVILEYE4 S_CPOS_DIE1 S_CPOS_DIE2 S_CPOS_DIE3 S_CPOS_DIE4 S_CPOS_DIE5 S_CPOS_DIE6 MAPBLOCKUNITS 128 HUSTR_E3M7 "E3M7: Limbo" S_CPOS_DIE7 mapped SPR_PLAS SIL_BOTTOM 1 AM_addMark GS_LEVEL __M_CONTROLS_H__  HUSTR_3 "level 3: the gantlet" S_TECH2LAMP S_BTORCHSHRT2 S_BSKULL2 key_flycenter ST_VERTICAL HUSTR_TALKTOSELF4 "You start to rave" SPR_PISG S_TBALL1 S_TBALL2 key_invhome dc_source S_BFGLAND2 S_BFGLAND3 S_BFGLAND4 S_BFGLAND5 S_BFGLAND6 deh_allow_long_strings S_SGUNUP PST_LIVE nodrawers transcolfunc SPR_TRE1 SPR_TRE2 key_lookcenter S_VILE_STND2 S_TECHLAMP4 ST_HEIGHT 32 MAXSWITCHES 50 SPR_TRED key_nextweapon S_PAIN_STND SCREENWIDTH_4_3 256 S_CPOS_STND2 S_PINS HUSTR_E2M7 "E2M7: Spawning Vats" S_PINV lastopening key_menu_qsave W_CacheLumpName exe_chex bfgedition amclock S_FATT_RAISE1 S_FATT_RAISE2 S_FATT_RAISE3 S_FATT_RAISE4 S_FATT_RAISE5 S_FATT_RAISE6 S_FATT_RAISE7 S_FATT_RAISE8 HUSTR_E1M1 "E1M1: Hangar" deathsound exe_hexen_1_1 ev_quit AM_drawMline key_spy key_arti_invulnerability AM_drawMarks video_driver tsilheight __P_LOCAL__  KEY_BACKSPACE 0x7f fastparm GAMMALVL2 "Gamma correction level 2" raiseAndChange __W_FILE__  S_CHAINFLASH1 S_CHAINFLASH2 key_strafeleft sk_hard tmpx HUSTR_E1M4 "E1M4: Command Control" am_noammo __AMMAP_H__  consistancy exe_heretic_1_3 it_bluecard HUSTR_11 "level 11: 'o' of destruction!" TSWALLRANGE GRAYSRANGE KEY_F1 (0x80+0x3b) S_SPOS_RAISE1 S_SPOS_RAISE2 S_SPOS_RAISE3 S_SPOS_RAISE4 ST_HORIZONTAL GOTSHELLS "Picked up 4 shotgun shells." AM_drawPlayers ML_BLOCKING 1 lowerToFloor joybmenu __P_PSPR__  key_menu_gamma AMSTR_FOLLOWOFF "Follow Mode OFF" parameter_chars key_invuse S_YSKULL2 weaponinfo S_CPOS_PAIN S_CSAW markpointnum key_menu_confirm levelTimeCount DOOUTCODE MAXINTERCEPTS_ORIGINAL 128 S_PAIN_ATK1 S_PAIN_ATK2 S_PAIN_ATK4 minx AM_maxOutWindowScale S_MEAT5 S_FATT_STND2 HUSTR_E1M8 "E1M8: Phobos Anomaly" S_PISTOLDOWN HUSTR_E2M2 "E2M2: Containment Area" KEY_F7 (0x80+0x41) LIGHTSCALESHIFT 12 blockbox S_SPOS_RAISE5 HUSTR_2 "level 2: underhalls" KEYP_PLUS '+' S_DSGUNFLASH2 netgame MT_WOLFSS S_PUNCH1 S_PUNCH2 S_PUNCH3 S_PUNCH4 S_PUNCH5 S_SPID_RUN3 S_SPID_RUN4 S_SPID_RUN5 S_SHOT2 S_SPID_RUN7 S_SPID_RUN8 S_SPID_RUN9 painsound NET_TICDIFF_CHATCHAR (1 << 5) key_arti_teleport S_TROO_STND2 wipegamestate exe_strife_1_2 MAXHEALTH 100 partime singledemo slopetype E1TEXT "Once you beat the big badasses and\n""clean out the moon base you're supposed\n""to win, aren't you? Aren't you? Where's\n""your fat reward and ticket home? What\n""the hell is this? It's not supposed to\n""end this way!\n""\n" "It stinks like rotten meat, but looks\n""like the lost Deimos base.  Looks like\n""you're stuck on The Shores of Hell.\n""The only way out is through.\n""\n""To continue the DOOM experience, play\n""The Shores of Hell and its amazing\n""sequel, Inferno!\n" playerstate HUSTR_E4M8 "E4M8: Unto The Cruel" SLOWDARK 35 __STSTUFF_H__  HUSTR_CHATMACRO4 "Help!" HUSTR_E4M4 "E4M4: Unruly Evil" S_BSPI_STND2 P5TEXT "You've found the second-hardest level we\n""got. Hope you have a saved game a level or\n""two previous.  If not, be prepared to die\n""aplenty. For master marines only." deathmatchstarts GOTBERSERK "Berserk!" thinglist doomstat.c dstrings.c EXIT_FAILURE 1 __INT_WCHAR_T_H  events RAND_MAX 0x7FFFFFFF _WCHAR_T_DEFINED_  result _BSD_WCHAR_T_ __WCHAR_T__  alloca __builtin_alloca __wchar_t__  MB_CUR_MAX 4 d_event.c __need_wchar_t __WCHAR_T  long long int __need_wchar_t  _WCHAR_T_DEFINED  D_PostEvent ___int_wchar_t_h  _T_WCHAR_  _WCHAR_T_DECLARED  _GCC_WCHAR_T  MLIBC_POSIX_STDLIB_H  _LOCALE_T_H  EXIT_SUCCESS 0 MLIBC_WCHAR_T_H  eventtail _T_WCHAR  D_PopEvent _BSD_WCHAR_T_  MAXEVENTS 64 eventhead _ALLOCA_H  d_items.c HAVE_LIBAMD64 IWAD_MASK_DOOM ((1 << doom) | (1 << doom2) | (1 << pack_tnt) | (1 << pack_plut) | (1 << pack_chex) | (1 << pack_hacx)) HAVE_LIBI386 SearchDirectoryForIWAD DirIsFile IWAD_MASK_HERETIC (1 << heretic) M_FileExists iwadfile strcasecmp d_iwad.c BuildIWADDirList iwad_dirs_built HAVE_LINUX_KD_H HAVE_DEV_ISA_SPKRIO_H PACKAGE "Doom" HAVE_LIBZ filename D_SaveGameIWADName M_StringJoin HAVE_SCHED_SETAFFINITY PACKAGE_TARNAME "doomgeneric.tar" iwads HAVE_LIBM iwad_t strcmp PACKAGE_STRING "Doom Generic 0.1" IdentifyIWADByName D_FindAllIWADs PACKAGE_VERSION 0.1 D_SuggestGameName num_iwad_dirs HAVE_MEMORY_H I_Error M_CheckParmWithArgs strrchr D_SuggestIWADName FILES_DIR "." D_FindIWAD _CTYPE_H  iwadname HAVE_LIBSAMPLERATE HAVE_MMAP HAVE_SYS_STAT_H PROGRAM_PREFIX "doomgeneric" HAVE_IOPERM MAX_IWAD_DIRS 128 CheckDirectoryHasIWAD STDC_HEADERS 1 HAVE_UNISTD_H __M_CONFIG__  PACKAGE_BUGREPORT configdir iwadparm HAVE_LIBPNG malloc strdup HAVE_DEV_SPEAKER_SPEAKER_H PACKAGE_NAME "Doom Generic" __D_IWAD__  IWAD_MASK_STRIFE (1 << strife) filename_len free IWAD_MASK_HEXEN (1 << hexen) D_TryFindWADByName result_len ORIGCODE AddIWADDir D_FindWADByName path_len d_loop.c SinglePlayerClear oldnettics FreeAddress num_players settings D_StartGameLoop AddrToString net_client_wait_data NET_SDL_H  BT_SPECIAL net_addr_t D_StartNetGame net_gamesettings_t ticcmd_set_t lasttime keyplayer _net_module_s players_mask availabletics gameticdiv _net_addr_s ticcmds NET_QUERY_H  net_server_wad_sha1sum net_broadcast_addr player_class I_Sleep nowtime net_packet_t BTS_SAVEMASK GetAdjustedTime RunMenu net_local_deh_sha1sum frameskip NET_IO_H  net_server_deh_sha1sum player_addrs recvtic RunTic NetUpdate BTS_PAUSE entertic net_local_is_freedoom SendPacket GetLowTic realtics net_server_is_freedoom net_connect_data_t new_sync BT_CHANGE ResolveAddress RecvPacket net_waiting_for_launch NET_SERVER_H  TicdupSquash _net_packet_s BTS_SAVEGAME BTS_SAVESHIFT respawn_monsters fast_monsters ready_players is_controller I_GetTime NET_GUI_H  NET_LOOP_H  skiptics newtics alloced D_InitNetGame net_module_t player_classes frameon BT_WEAPONSHIFT ticdata net_sdl_module net_loop_client_module I_StartTic net_local_wad_sha1sum D_RegisterLoopCallbacks I_AtExit maketic NET_CLIENT_H  net_waitdata_t oldentertics max_players connect_data D_ReceiveTic BuildNewTic extratics InitServer TryRunTics net_client_received_wait_data local_playeringame BT_ATTACK net_loop_server_module num_drones player_names PlayersInGame OldNetSync offsetms random loop_interface_t BT_WEAPONMASK I_GetTimeMS D_QuitNetGame localplayer sha1_digest_t handle InitClient lowtic BT_USE BT_SPECIALMASK netgame_startup_callback_t net_player_name D_Disconnected I_SetWindowTitle HU_BROADCAST 5 __P_SETUP__  link I_BindJoystickVariables D_BindVariables __P_SAVEG__  mus_romer2 snd_maxslicetime_ms W_MAIN_H  HU_MSGWIDTH 64 D_AdvanceDemo driver_data gameversions advancedemo I_PrintStartupBanner __M_MENU__  viewactivestate HU_FONTSIZE (HU_FONTEND - HU_FONTSTART + 1) G_InitNew M_BindChatControls sfxinfo_t snd_musicdevice R_Init sfxinfo_struct R_DrawViewBorder W_CheckNumForName ga_newgame HAT_AXIS_HORIZONTAL 1 D_IdentifyVersion I_InitSound M_LoadDefaults mus_romero mus_count2 atoi InitGameVersion gameaction mus_countd wipe_NUMWIPES ST_Drawer I_DisplayFPSDots V_Init IS_BUTTON_AXIS(axis) ((axis) >= 0 && ((axis) & BUTTON_AXIS) != 0) I_InitGraphics V_DrawPatchDirect demosequence deh_sub HU_FONTSTART '!' mus_dead2 gameaction_t HU_FONTEND '_' W_AddFile NUMMUSIC snd_cachesize mus_dm2int I_FinishUpdate SetMissionForPackName mus_e2m1 mus_e2m2 mus_e2m3 mus_e2m4 mus_e2m5 mus_e2m6 mus_e2m7 mus_e2m8 mus_e2m9 M_BindVariable wipe_ColorXForm G_TimeDemo I_StartFrame strncasecmp is_freedm ga_loadlevel tagname D_StartTitle __I_JOYSTICK__  M_StringCopy SAVESTRINGSIZE 24 mus_read_m vanilla_demo_limit I_PrintBanner mus_stlks3 mus_dm2ttl HU_MSGY 0 I_InitJoystick demolumpname V_RestoreBuffer wipestart I_BindVideoVariables I_SetPalette numchannels mus_introa __WI_STUFF__  deh_s W_CheckCorrectIWAD D_CheckNetGame I_PrintDivider showMessages ga_loadgame wipe_Melt HAT_AXIS_VERTICAL 2 storedemo oldgamestate screenblocks __F_WIPE_H__  G_Responder V_DrawMouseSpeedBox borderdrawcount mus_stalks mus_dead I_InitMusic M_StringEndsWith R_ExecuteSetViewSize usefulness save_stream NET_DEDICATED_H  mus_betwee mapdir M_BindBaseControls mus_ddtbl2 mus_ddtbl3 mus_ddtblu atexit_func_t S_Init snd_musiccmd wipe_ScreenWipe mus_theda2 mus_theda3 ga_playdemo I_UpdateNoBlit W_ParseCommandLine DOOM_STATDUMP_H  D_AddFile D_Endoom M_BindMapControls M_BindMenuControls mus_openin G_BeginRecording S_sfx gamename_size mus_evil mus_e3m2 mus_victor I_CheckIsScreensaver P_Init copyright_banners vanilla_savegame_limit R_FillBackScreen CREATE_BUTTON_AXIS(neg,pos) (BUTTON_AXIS | (neg) | ((pos) << 8)) HAT_AXIS_DIRECTION(axis) (((axis) >> 8) & 0xff) ST_Init I_InitTimer pagetic D_ConnectNetGame F_Drawer ga_worlddone M_Init G_RecordDemo HU_Init M_SetConfigFilenames BUTTON_AXIS_POS(axis) (((axis) >> 8) & 0xff) mus_shawn2 mus_shawn3 D_DoomLoop CREATE_HAT_AXIS(hat,direction) (HAT_AXIS | (hat) | ((direction) << 8)) inhelpscreensstate pagename mus_bunny HAT_AXIS_HAT(axis) ((axis) & 0xff) G_LoadGame setsizeneeded Z_Init HU_MSGTIMEOUT (4*TICRATE) __S_SOUND__  NUM_VIRTUAL_BUTTONS 10 wipe_StartScreen GetGameName ga_savegame mus_runni2 musicinfo_t snd_sfxdevice packs gamename menuactivestate M_BindWeaponControls __G_GAME__  __F_FINALE__  ga_victory BUTTON_AXIS_NEG(axis) ((axis) & 0xff) HU_MSGHEIGHT 1 mus_runnin S_UpdateSounds mus_e1m1 mus_e1m2 mus_e1m3 mus_e1m4 mus_e1m5 mus_e1m6 mus_e1m7 mus_e1m8 mus_e1m9 HU_MSGX 0 __SOUNDS__  d_main.c ga_completed HAT_AXIS 0x20000 chat_macros HU_Erase M_ApplyPlatformDefaults mus_adrian I_EnableLoadingDisk __I_SOUND__  show_endoom main_loop_started mus_ampie ga_screenshot savegame_error I_SetGrabMouseCallback PrintDehackedBanners WI_Drawer D_GrabMouseCallback redrawsbar mus_e3m1 mus_e3m3 mus_e3m4 mus_e3m5 mus_e3m6 mus_e3m7 mus_e3m8 mus_e3m9 S_music mus_stlks2 M_CheckParm mus_ultima __D_MAIN__  pack_name D_Display __HU_STUFF_H__  I_BindSoundVariables mus_shawn D_ProcessEvents detailLevel M_GetSaveGameDir mus_inter PrintGameVersion mus_None mus_messag __I_ENDOOM__  D_PageTicker ga_nothing D_PageDrawer mus_doom2 mus_tense I_Endoom mus_messg2 snd_samplerate D_DoAdvanceDemo wipe inhelpscreens snd_channels G_DeferedPlayDemo mus_in_cit D_SetGameDescription W_GenerateHashTable S_StartMusic IS_HAT_AXIS(axis) ((axis) >= 0 && ((axis) & HAT_AXIS) != 0) HU_Drawer cmdline mus_intro M_SetConfigDir mus_doom R_RenderPlayerView P_SaveGameFile I_GraphicsCheckCommandLine BUTTON_AXIS 0x10000 mus_the_da wipe_EndScreen D_IsEpisodeMap valid_modes D_ValidGameMode D_GetNumEpisodes D_ValidEpisodeMap d_mode.c valid_versions D_ValidGameVersion D_GameMissionString player_num W_Checksum LoadGameSettings G_CheckDemoStatus exitmsg W_CHECKSUM_H  doom_loop_interface SaveGameSettings PlayerQuitGame InitConnectData G_Ticker d_net.c __builtin_putchar sfx_popain F_STAGE_ARTSCREEN sfx_posit1 sfx_posit3 sfx_sklatk sfx_sawhit sfx_sawful sfx_plasma sfx_bossit f_finale.c sfx_radio castnum sfx_sgtatk sfx_stnmov sfx_pistol sfx_dbcls NUMSFX F_BunnyScroll sfx_pedth sfx_bgdth2 event F_ArtScreenDrawer sfx_podth1 sfx_podth2 sfx_podth3 F_TextWrite sprframe sfx_spidth sfx_getpow S_StartSound sfx_itmbk textscreen_t sfx_skedth sfx_bgact sfx_dorcls V_DrawPatchFlipped sfx_bdcls sfx_ssdth hu_font S_ChangeMusic casttics sfx_kntdth sfx_noway sfx_mnpain castdeath sfx_spisit toupper post_t scrolled sfx_vilsit sfx_dmpain sfx_vipain F_STAGE_TEXT W_CacheLumpNum topdelta finaletext sfx_sssit __I_SWAP__  sfx_boscub sfx_bspdth sfx_sgcock TEXTSPEED 3 sfx_dbload sfx_brsdth sfx_wpnup F_CastDrawer caststate sfx_bospit sfx_bgsit1 sfx_bgsit2 sfx_kntsit sfx_oof sfx_cacdth F_CastPrint TEXTWAIT 250 desttop sfx_keendt sfx_telept sfx_rxplod SHORT(x) ((signed short) (x)) sfx_flame sfx_pstop sfx_bosdth F_STAGE_CAST sfx_posact F_Responder LONG(x) ((signed int) (x)) sfx_bspsit sfx_brssit sfx_chgun sfx_swtchx sfx_pesit sfx_swtchn sfx_vilact F_StartCast textscreens F_DrawPatchCol sfx_cybdth sfx_punch sfx_sawidl sfx_vilatk sfx_skldth sfx_keenpn stopattack sfx_pldeth sfx_bspact sfx_hoof background sfx_slop sfx_mandth sfx_barexp F_StartFinale sfx_None sfx_firsht castinfo_t sfx_itemup finalestage_t sfx_tink sfx_skesit sfx_cybsit castframes sfx_bfg sfx_flamst F_CastResponder sfx_dbopn sfx_cacsit sfx_sgtdth sfx_sawup sfx_bspwlk column_t sfx_mansit sfx_bgdth1 sfx_skeact sfx_rlaunc sfx_skeswg sfx_doropn sfx_dmact sfx_sgtsit sfx_firxpl sfx_pdiehi sfx_pepain sfx_metal F_CastTicker castorder sprdef castonmelee sfx_skeatk sfx_dshtgn sfx_bospn sfx_shotgn castattacking finaleflat laststage sfx_manatk sfx_bdopn sfx_pstart finalecount sfx_plpain sfx_posit2 sfx_vildth sfx_skepch SYS_LITTLE_ENDIAN  sfx_claw finalestage F_Ticker Z_Free wipe_doColorXForm wipe_scr newval changed wipeno I_ReadScreen __M_RANDOM__  V_DrawBlock wipe_scr_start wipes ticks wipe_doMelt f_wipe.c wipe_shittyColMajorXform wipe_exitMelt wipe_initColorXForm wipe_initMelt M_Random wipe_scr_end wipe_exitColorXForm Z_Malloc P_ArchiveSpecials new_length dclickstate2 _MATH_H  __R_SKY__  netdemo P_WriteSaveGameEOF isless(x,y) __MLIBC_CHOOSE_COMPARISON(x, y, __mlibc_isless) DEH_DEFAULT_SPECIES_INFIGHTING 0 P_Random buttons_mask DEH_DEFAULT_BLUE_ARMOR_CLASS 2 WI_Ticker G_ReadDemoTiccmd M_LOG2E 1.4426950408889634074 P_SpawnPlayer turbodetected d_skill MF_TELEPORT IncreaseDemoBuffer P_WriteSaveGameHeader Z_CheckHeap DEH_DEFAULT_GOD_MODE_HEALTH 100 __P_TICK__  joyymove M_LOG10E 0.43429448190325182765 savegameslot deh_idfa_armor DEH_DEFAULT_IDFA_ARMOR G_DeferedInitNew M_2_SQRTPI 1.12837916709551257390 P_ArchivePlayers V_ScreenShot DEH_DEFAULT_IDKFA_ARMOR_CLASS 2 DEH_DEFAULT_MAX_SOULSPHERE 200 DEH_DEFAULT_INITIAL_HEALTH 100 savedleveltime temp_savegame_file M_1_PI 0.31830988618379067154 FP_ILOGBNAN (-1 - (int)(((unsigned)-1) >> 1)) TURBOTHRESHOLD 0x32 turbomessage G_DoNewGame new_demop g_game.c MAX_JOY_BUTTONS 20 skytexturemid savedescription DEH_DEFAULT_IDFA_ARMOR_CLASS 2 MAXPLMOVE (forwardmove[1]) ANGLETOSKYSHIFT 22 M_StartControlPanel turnheld signbit(x) (__builtin_signbit(x)) MF_TRANSSHIFT G_PlayerFinishLevel MF_SHOOTABLE P_SetupLevel secretexit sendpause M_LN2 0.69314718055994530942 R_TextureNumForName BODYQUESIZE 32 MF_SPECIAL deh_max_armor DEH_DEFAULT_MAX_ARMOR G_CheckSpot DEH_DEFAULT_GREEN_ARMOR_CLASS 1 MF_JUSTATTACKED M_SQRT2 1.41421356237309504880 S_PauseSound dclicktime MF_SKULLFLY M_SQRT1_2 0.70710678118654752440 HUGE_VAL (__builtin_huge_val()) mousex mousey FP_ZERO 16 P_CheckPosition weapon_keys button_on G_NextWeapon MF_SPAWNCEILING MF_MISSILE sendsave HUGE_VALL (__builtin_huge_vall()) playernum MF_NOBLOCKMAP G_BuildTiccmd dclicks isinf(x) (fpclassify(x) == FP_INFINITE) cpars MF_NOGRAVITY demoversion G_SecretExitLevel SetJoyButtons isnan(x) (fpclassify(x) == FP_NAN) M_PI_4 0.78539816339744830962 resultbuf demoname_size MF_DROPOFF joybuttons DEH_DEFAULT_MAX_ARMOR 200 DEH_DEFAULT_MEGASPHERE_HEALTH 200 HU_Ticker ST_Ticker deh_initial_health DEH_DEFAULT_INITIAL_HEALTH G_SaveGame MF_INFLOAT joyarray M_LN10 2.30258509299404568402 WI_Start bodyque P_ReadSaveGameEOF FP_INFINITE 1 dclicktime2 MF_COUNTITEM NUMKEYS 256 NAN (__builtin_nanf("")) d_episode MF_NOCLIP desired_angleturn defdemoname islessgreater(x,y) __MLIBC_CHOOSE_COMPARISON(x, y, __mlibc_islessgreater) deh_max_health DEH_DEFAULT_MAX_HEALTH G_DeathMatchSpawnPlayer S_ResumeSound dclicks2 DEH_DEFAULT_INITIAL_BULLETS 50 MF_SOLID MF_JUSTHIT deh_green_armor_class DEH_DEFAULT_GREEN_ARMOR_CLASS SKYFLATNAME "F_SKY1" joystrafemove P_ReadSaveGameHeader starttime start_i current_length deh_blue_armor_class DEH_DEFAULT_BLUE_ARMOR_CLASS demo_start DemoVersionDescription remove MF_TRANSLATION G_DoPlayDemo G_VanillaVersionCode weapon_order_table P_UnArchivePlayers maxsize FP_NORMAL 4 selections G_DoWorldDone MATH_ERREXCEPT 2 deh_bfg_cells_per_shot DEH_DEFAULT_BFG_CELLS_PER_SHOT P_ArchiveThinkers deh_species_infighting DEH_DEFAULT_SPECIES_INFIGHTING deh_max_soulsphere DEH_DEFAULT_MAX_SOULSPHERE MF_NOSECTOR M_ClearRandom DEMOMARKER 0x80 recovery_savegame_file P_SpawnMobj P_ArchiveWorld isunordered(x,y) (isnan((x)) ? ((void)(y),1) : isnan((y))) R_FlatNumForName M_PI_2 1.57079632679489661923 isgreater(x,y) __MLIBC_CHOOSE_COMPARISON(x, y, __mlibc_isgreater) mousebuttons skytexturename P_UnArchiveWorld G_WorldDone FP_NAN 2 WI_End MF_SLIDE deh_idkfa_armor_class DEH_DEFAULT_IDKFA_ARMOR_CLASS VERSIONSIZE 16 deh_idkfa_armor DEH_DEFAULT_IDKFA_ARMOR M_PI 3.14159265358979323846 savename G_CmdChecksum isfinite(x) (fpclassify(x) & (FP_NORMAL | FP_SUBNORMAL | FP_ZERO)) __MLIBC_CHOOSE_COMPARISON(x,y,p) ( sizeof((x)+(y)) == sizeof(float) ? p ##f(x, y) : sizeof((x)+(y)) == sizeof(double) ? p(x, y) : p ##l(x, y) ) deh_god_mode_health DEH_DEFAULT_GOD_MODE_HEALTH G_DoCompleted demoend fpclassify(x) (sizeof(x) == sizeof(double) ? __fpclassify(x) : (sizeof(x) == sizeof(float) ? __fpclassifyf(x) : (sizeof(x) == sizeof(long double) ? __fpclassifyl(x) : 0))) R_PointInSubsector deh_idfa_armor_class DEH_DEFAULT_IDFA_ARMOR_CLASS FP_SUBNORMAL 8 DEH_DEFAULT_BFG_CELLS_PER_SHOT 40 DEH_DEFAULT_MAX_HEALTH 200 carry P_Ticker d_map G_DoSaveGame isnormal(x) (fpclassify(x) == FP_NORMAL) skytexture G_InitPlayer timingdemo dclickstate weapon_num next_weapon MF_NOTDMATCH MF_NOBLOOD StatCopy islessequal(x,y) __MLIBC_CHOOSE_COMPARISON(x, y, __mlibc_islessequal) G_PlayerReborn MF_PICKUP SetMouseButtons endtime M_E 2.7182818284590452354 G_DoLoadLevel HUGE_VALF (__builtin_huge_valf()) P_UnArchiveThinkers M_2_PI 0.63661977236758134308 deh_megasphere_health DEH_DEFAULT_MEGASPHERE_HEALTH INFINITY (__builtin_inff()) G_ExitLevel MF_CORPSE tspeed HU_dequeueChatChar WeaponSelectable M_WriteFile MF_COUNTKILL I_Quit deh_initial_bullets DEH_DEFAULT_INITIAL_BULLETS mousearray FP_ILOGB0 FP_ILOGBNAN DEH_MISC_H  joyxmove fopen G_ScreenShot P_TempSaveGameFile G_DoLoadGame DEH_DEFAULT_SOULSPHERE_HEALTH 100 math_errhandling 3 P_UnArchiveSpecials G_WriteDemoTiccmd MF_AMBUSH MF_FLOAT MF_DROPPED HU_Responder deh_soulsphere_health DEH_DEFAULT_SOULSPHERE_HEALTH MF_SHADOW new_demobuffer DEH_DEFAULT_IDFA_ARMOR 200 isgreaterequal(x,y) __MLIBC_CHOOSE_COMPARISON(x, y, __mlibc_isgreaterequal) DEH_DEFAULT_IDKFA_ARMOR 200 longtics MATH_ERRNO 1 G_DoReborn demo_p P_RemoveMobj M_TempFile SLOWTURNTICS 6 SAVEGAMESIZE 0x2c000 gamekeydown drawcursor needsupdate R_VideoErase HUlib_drawTextLine HUlib_delCharFromIText hu_textline_t HUlib_keyInIText startchar HUlib_drawIText HUlib_delCharFromTextLine hu_itext_t HUlib_addCharToTextLine HUlib_initIText HU_CHARERASE KEY_BACKSPACE __HULIB__  HUlib_clearTextLine HUlib_eraseIText yoffset hu_stext_t HUlib_addLineToSText HUlib_addMessageToSText HUlib_eraseSText HUlib_initSText HUlib_drawSText HUlib_addPrefixToIText HUlib_initTextLine HUlib_init HUlib_eraseTextLine laston HU_MAXLINES 4 HUlib_resetIText noterased viewwindowx hu_lib.c HUlib_eraseLineFromIText HU_MAXLINELENGTH 80 HU_Stop HU_TITLE (mapnames[(gameepisode-1)*9+gamemap-1]) HU_TITLEHEIGHT 1 HU_INPUTWIDTH 64 HU_INPUTY (HU_MSGY + HU_MSGHEIGHT*(SHORT(hu_font[0]->height) +1)) HU_TITLE_CHEX (mapnames[gamemap - 1]) w_title HU_queueChatChar mapnames_commercial chat_char HU_Start QUEUESIZE 128 message_on HU_TITLEY (167 - SHORT(hu_font[0]->height)) altdown num_nobrainers headsupactive message_counter message_nottobefuckedwith chat_dest w_chat eatkey always_off HU_TITLET (mapnames_commercial[gamemap-1 + 64]) message_dontfuckwithme mapnames chatchars w_inputbuffer chat_on numplayers HU_TITLEP (mapnames_commercial[gamemap-1 + 32]) HU_TITLEX 0 macromessage HU_INPUTX HU_MSGX HU_TITLE2 (mapnames_commercial[gamemap-1]) HU_INPUTTOGGLE 't' HU_INPUTHEIGHT 1 lastmessage hu_stuff.c w_message info.c __ICDMUS__  CDERR_DEVREQBASE 100 cd_Error track CDERR_NOTINSTALLED 10 I_CDMusInit I_CDMusPrintStartup CDERR_BADTRACK 21 CDERR_IOCTLBUFFMEM 22 I_CDMusTrackLength I_CDMusResume I_CDMusSetVolume I_CDMusFirstTrack I_CDMusStop track_num CDERR_NOAUDIOSUPPORT 11 CDERR_BADDRIVE 20 I_CDMusPlay i_cdmus.c CDERR_NOAUDIOTRACKS 12 I_CDMusLastTrack endoom_data ENDOOM_W 80 ENDOOM_H 25 i_endoom.c usejoystick I_ShutdownJoystick joystick_strafe_axis joystick_physical_buttons joystick_x_axis joystick_y_invert joystick_y_axis joystick_index joystick_x_invert joystick_strafe_invert i_joystick.c DEAD_ZONE (32768 / 3) I_UpdateJoystick col1 I_InitSquashTable dest2 dest3 dest4 dest5 screenp I_ResetScaleTables col2 I_Scale2x I_Scale5x DrawScreen WriteSquashedLine1x I_Scale1x WriteSquashedLine2x i_scale.c WriteSquashedLine3x multi_pitch I_InitScale mode_scale_1x WriteLine3x InitMode WriteSquashedLine5x _dest_pitch mode_scale_2x mode_scale_5x mode_scale_3x _dest_buffer I_InitStretchTables mode_scale_4x WriteBlendedLine1x I_Squash1x WriteBlendedLine2x mode_squash_1x I_Squash2x bufp WriteLine2x I_Squash3x mode_squash_2x WriteBlendedLine4x I_Squash4x mode_squash_3x mode_stretch_1x WriteLine4x I_Squash5x mode_squash_4x mode_stretch_4x mode_stretch_2x WriteLine5x mode_squash_5x mode_stretch_3x I_Stretch1x screenp4 src2 I_Stretch2x src1 FindNearestColor mode_stretch_5x best GenerateStretchTable I_Stretch3x half_stretch_table I_Stretch4x screen_mode_t I_Stretch5x I_Scale3x WriteSquashedLine4x _src_buffer WriteBlendedLine3x I_Scale4x best_diff DRAW_PIXEL2 *dest++ = *dest2++ = c; DRAW_PIXEL4 *dest++ = *dest2++ = *dest3++ = *dest4++ = c; stretch_tables DRAW_PIXEL5 *dest++ = *dest2++ = *dest3++ = *dest4++ = *dest5++ = c DRAW_PIXEL3 *dest++ = *dest2++ = *dest3++ = c fflush screenp2 screenp3 poor_quality screenp5 I_PrecacheSounds music_opl_module SndDeviceInList sound_sdl_module CheckVolumeSeparation nomusic I_StopSound PauseMusic SNDDEVICE_PCSPEAKER I_SetMusicVolume CacheSounds InitSfxModule nosfx timidity_cfg_path num_sounds music_module num_sound_devices I_MusicIsPlaying I_StopSong SNDDEVICE_ADLIB use_sfx_prefix I_SoundIsPlaying looping I_PlaySong I_UnRegisterSong I_UpdateSound I_PauseSong I_ShutdownMusic SNDDEVICE_SB channel SNDDEVICE_GUS SNDDEVICE_AWE32 music_modules SNDDEVICE_NONE I_StartSound I_ResumeSong I_RegisterSong SNDDEVICE_PAS SNDDEVICE_WAVEBLASTER opl_io_port I_ShutdownSound nosound InitMusicModule i_sound.c SNDDEVICE_SOUNDCANVAS ResumeMusic music_module_t sound_module_t sound_pcsound_module Poll I_GetSfxLumpNum SNDDEVICE_CD I_UpdateSoundParams sfxinfo music_sdl_module sound_modules snddevice_t SNDDEVICE_GENMIDI ZenityErrorBox _CS_POSIX_V6_ILP32_OFFBIG_LIBS 1122 errorboxpath_size _CS_POSIX_V6_ILP32_OFFBIG_LINTFLAGS 1123 ZENITY_BINARY "/usr/bin/zenity" _PC_NAME_MAX 3 _CS_PATH 0 _CS_POSIX_V5_WIDTH_RESTRICTED_ENVS 4 _CS_GNU_LIBPTHREAD_VERSION 3 spaces zonemem STDIN_FILENO 0 mem_dump_win98 STDOUT_FILENO 1 _CS_POSIX_V6_ILP32_OFFBIG_LDFLAGS 1121 _SC_OPEN_MAX 5 _SC_PAGE_SIZE 3 MIN_RAM 6 _CS_POSIX_V7_ILP32_OFFBIG_LINTFLAGS 1139 _CS_POSIX_V6_LP64_OFF64_CFLAGS 1124 dos_mem_dump _CS_POSIX_V7_ILP32_OFF32_CFLAGS 1132 _UNISTD_H  system environ _CS_POSIX_V6_WIDTH_RESTRICTED_ENVS 1 _CS_POSIX_V6_LP64_OFF64_LDFLAGS 1125 __gnuc_va_list F_OK 1 _CS_POSIX_V7_ILP32_OFF32_LDFLAGS 1133 ZenityAvailable I_ZoneBase X_OK 8 exit_gui_popup run_on_error _CS_POSIX_V7_ILP32_OFFBIG_CFLAGS 1136 F_TLOCK 3 W_OK 4 __va_list_tag _CS_POSIX_V6_ILP32_OFF32_LINTFLAGS 1119 _CS_POSIX_V6_LPBIG_OFFBIG_LIBS 1130 _SC_ARG_MAX 0 I_Tactile MLIBC_GID_T_H  optind _CS_POSIX_V7_ILP32_OFFBIG_LDFLAGS 1137 _CS_POSIX_V7_WIDTH_RESTRICTED_ENVS 5 exit_funcs _CS_POSIX_V7_ILP32_OFF32_LINTFLAGS 1135 errorboxpath reg_save_area _PC_LINK_MAX 0 i_system.c _CS_POSIX_V6_LPBIG_OFFBIG_LDFLAGS 1129 F_ULOCK 4 F_LOCK 1 mem_dump_dosbox __builtin_fputs __builtin_va_list gp_offset DOS_MEM_DUMP_SIZE 10 _CS_POSIX_V7_ILP32_OFF32_LIBS 1134 _PC_PATH_MAX 4 overflow_arg_area MLIBC_PID_T_H  total AutoAllocMemory _CS_POSIX_V7_ILP32_OFFBIG_LIBS 1138 _SC_GETPW_R_SIZE_MAX 1 msgbuf atexit_listentry_s atexit_listentry_t _CS_POSIX_V6_LPBIG_OFFBIG_LINTFLAGS 1131 M_vsnprintf _CS_POSIX_V7_LPBIG_OFFBIG_CFLAGS 1144 already_quitting entry DEFAULT_RAM 6 optopt mem_dump_custom _CS_POSIX_V6_ILP32_OFF32_LDFLAGS 1117 escaped_message _CS_POSIX_V6_LP64_OFF64_LIBS 1126 mem_dump_dos622 opterr _CS_POSIX_V6_ILP32_OFF32_LIBS 1118 fp_offset _CS_V7_ENV 1149 _XOPEN_VERSION 700 _CS_POSIX_V6_LPBIG_OFFBIG_CFLAGS 1128 _CS_POSIX_V7_LPBIG_OFFBIG_LDFLAGS 1145 strchr I_ConsoleStdout default_ram _CS_POSIX_V7_LP64_OFF64_LDFLAGS 1141 _SC_PAGESIZE _SC_PAGE_SIZE _CS_V6_ENV 1148 I_GetMemoryValue _CS_GNU_LIBC_VERSION 2 _CS_POSIX_V7_LP64_OFF64_CFLAGS 1140 _CS_POSIX_V7_LPBIG_OFFBIG_LINTFLAGS 1147 F_TEST 2 _POSIX2_VERSION 200809L _SC_PHYS_PAGES 2 _CS_POSIX_V7_LP64_OFF64_LIBS 1142 STDERR_FILENO 2 _CS_POSIX_V7_LP64_OFF64_LINTFLAGS 1143 _PC_PIPE_BUF 5 _CS_POSIX_V6_LP64_OFF64_LINTFLAGS 1127 _POSIX_THREADS 200809L argptr _POSIX_VERSION 200809L optarg M_ParmExists R_OK 2 M_StrToInt min_ram _CS_POSIX_V7_LPBIG_OFFBIG_LIBS 1146 MLIBC_UID_T_H  _CS_POSIX_V6_ILP32_OFFBIG_CFLAGS 1120 EscapeShellString _CS_POSIX_V6_ILP32_OFF32_CFLAGS 1116 vfprintf __mlibc_uint32 uint32_t basetime DOOMGENERIC_RESY 400 DOOMGENERIC_RESX 640 DG_SleepMs DG_ScreenBuffer DOOM_GENERIC  I_WaitVBL DG_GetTicksMs I_GetTicks i_timer.c mem_rel_t mem_fread MEM_SEEK_CUR newbuf memio.c mem_get_buf _MEMFILE newpos MODE_READ MEMIO_H  MEM_SEEK_SET buflen MEM_SEEK_END MODE_WRITE nmemb mem_fclose whence memfile_mode_t mem_fseek mem_fopen_write mem_ftell mem_fopen_read mem_fwrite LoadResponseFile MAXARGVS 100 m_argv.c M_GetExecutableName num_args argv_index M_ClearBox M_AddToBox BOXTOP BOXRIGHT BOXLEFT BOXBOTTOM __M_BBOX__  m_bbox.c cht_GetParam m_cheat.c ENFILE 1040 EINPROGRESS 1024 EPROTO 1065 ECONNREFUSED 1014 DEFAULT_INT M_SetVariable ENOTCONN 1052 EINTR 1025 doom_defaults_list ENOENT 1043 EFAULT 1020 atof original_translated ECANCELED 1011 ETXTBSY 1073 GetDefaultForName M_GetStrVariable ENOTRECOVERABLE 1055 ENOTSUP 1057 default_type_t DEFAULT_KEY EBUSY 1010 CONFIG_VARIABLE_GENERIC(name,type) { #name, NULL, type, 0, 0, false } EDEADLK 1016 EOPNOTSUPP 1060 EBADMSG 1009 CONFIG_VARIABLE_KEY(name) CONFIG_VARIABLE_GENERIC(name, DEFAULT_KEY) ENETRESET 1038 ENODEV 1042 EOVERFLOW 1061 ENXIO 1059 ERANGE 3 errno __mlibc_errno EMFILE 1031 ENOEXEC 1044 ESPIPE 1069 ENOPROTOOPT 1049 EISDIR 1029 ENOKEY 1078 ENOTDIR 1053 LoadDefaultCollection EACCES 1002 DEFAULT_INT_HEX ELOOP 1030 orig_extra EHOSTUNREACH 1022 ENOTTY 1058 E2BIG 1001 default_t program_invocation_name SaveDefaultCollection ENOSPC 1050 ENOBUFS 1041 CONFIG_VARIABLE_INT(name) CONFIG_VARIABLE_GENERIC(name, DEFAULT_INT) ENODATA 1076 default_collection_t strparm ENETUNREACH 1039 ETIMEDOUT 1072 EDQUOT 1018 location _ABIBITS_ERRNO_H  ENOMSG 1048 EDESTADDRREQ 1017 intparm M_SaveDefaults EPERM 1063 ENOLCK 1045 EALREADY 1007 scantokey sscanf EADDRNOTAVAIL 1004 EADDRINUSE 1003 ETIME 1077 ENAMETOOLONG 1036 m_config.c EIDRM 1023 DEFAULT_FLOAT ESTALE 1071 EBADF 1008 EXDEV 1075 default_main_config orig_main CONFIG_VARIABLE_INT_HEX(name) CONFIG_VARIABLE_GENERIC(name, DEFAULT_INT_HEX) ENOSYS 1051 EMSGSIZE 1034 variable EINVAL 1026 ParseIntParameter M_GetFloatVariable CONFIG_VARIABLE_STRING(name) CONFIG_VARIABLE_GENERIC(name, DEFAULT_STRING) extra_defaults_list bound program_invocation_short_name ESRCH 1070 EPROTOTYPE 1067 ECHILD 1012 EEXIST 1019 EAGAIN 1006 SearchCollection EPIPE 1064 EROFS 1068 EPROTONOSUPPORT 1066 extra_defaults ENOMEM 1047 EOWNERDEAD 1062 CONFIG_VARIABLE_FLOAT(name) CONFIG_VARIABLE_GENERIC(name, DEFAULT_FLOAT) M_MakeDirectory numdefaults DEFAULT_STRING ENETDOWN 1037 GetDefaultConfigDir M_SaveDefaultsAlternate EAFNOSUPPORT 1005 EFBIG 1021 doom_defaults EILSEQ 2 EMULTIHOP 1035 default_extra_config EDOM 1 ENOTSOCK 1056 M_GetIntVariable EWOULDBLOCK EAGAIN ECONNABORTED 1013 EIO 1027 ECONNRESET 1015 untranslated EMLINK 1032 collection EISCONN 1028 ENOLINK 1046 ENOTEMPTY 1054 M_BindStrifeControls m_controls.c M_BindHexenControls M_BindHereticControls __mlibc_int64 m_fixed.c newg_end M_DrawSelCell M_DoSave currentMenu quitsounds read1_end M_DrawSound M_DrawEpisode rdthsempty2 gammamsg messageNeedsInput M_ReadSaveStrings mousesens SaveMenu M_SaveSelect EpiDef hurtme M_SaveGame killthings messageRoutine quitdoom skullAnimCounter M_FinishReadThis sfx_empty1 prevMenu toorough M_QuickLoadResponse IsNullKey M_EndGame option_empty2 sfx_vol quitsounds2 itemOn violence M_ChangeDetail M_QuitResponse SKULLXOFF -32 choice M_LoadGame detailNames M_ChangeMessages OptionsMenu M_DrawThermo load_e M_StringWidth M_QuickLoad read_e2 sound_e saveStringEnter tempstring M_DrawReadThis1 M_DrawReadThis2 S_SetMusicVolume option_empty1 music_vol msgNames input messageString thermDot sound_end readthis episodes_e saveCharIndex SoundMenu whichSkull NewGameMenu M_DrawSave ReadDef1 ReadDef2 read2_end sfx_empty2 quickSaveSlot LoadMenu skullName ep_end thermWidth M_NewGame M_Options M_MusicVol M_ChangeSensitivity M_Sound ReadMenu1 ReadMenu2 SoundDef M_StringHeight load_end savegamestrings options_e foundnewline routine M_QuickSaveResponse M_ChooseSkill M_ClearMenus screenSize M_VerifyNightmare joywait read_e M_DrawSaveLoadBorder scrnsize M_SelectEndMessage mousewait M_StopMessage main_e saveSlot rdthsempty1 main_end opt_end M_StartMessage newgame_e EpisodeMenu LINEHEIGHT 16 menudef endstring menu_s menu_t skullx skully menuitem_t item M_SfxVol M_DrawNewGame M_DrawOptions M_ReadThis2 saveOldString m_menu.c M_SetupNextMenu M_WriteText R_SetViewSize lastOn M_Episode M_EndGameResponse messageToPrint lastx lasty S_SetSfxVolume M_QuitDOOM load1 load4 load6 messx messy M_LoadSelect M_DrawEmptyCell soundvol OptionsDef menuitems messageLastMenuActive numitems M_QuickSave alphaKey load2 load3 load5 MainDef SaveDef M_SizeDisplay M_DrawLoad LoadDef M_ReadThis NewDef M_DrawMainMenu replacement st_atime st_atim.tv_sec M_StringReplace MLIBC_MODE_T_H  S_IXGRP 010 S_IFCHR 0x02000 M_FileLength S_IWOTH 02 _ABIBITS_STAT_H  MLIBC_TIME_T  MLIBC_NLINK_T_H  MLIBC_BLKCNT_T_H  dst_len S_ISVTX 01000 MLIBC_STAT_H  MLIBC_FSBLKCNT_T_H  _SYS_TYPES_H  MLIBC_FSFILCNT_T_H  st_mtime st_mtim.tv_sec S_IROTH 04 m_misc.c S_IRWXU 0700 mkdir S_IRGRP 040 S_IRWXO 07 S_IWUSR 0200 haystack_len S_IXUSR 0100 M_ExtractFileBase S_ISREG(m) (((m) & S_IFMT) == S_IFREG) S_IWGRP 020 needle S_ISLNK(m) (((m) & S_IFMT) == S_IFLNK) S_ISSOCK(m) (((m) & S_IFMT) == S_IFSOCK) fstream S_ISGID 02000 S_ISDIR(m) (((m) & S_IFMT) == S_IFDIR) S_IFSOCK 0x0C000 S_IFLNK 0x0A000 M_ReadFile savedpos dest_size needle_len M_StringConcat orig suffix S_ISUID 04000 strncmp S_IRWXG 070 S_IFBLK 0x06000 MLIBC_SUSECONDS_T_H  tempdir st_ctime st_ctim.tv_sec S_IFMT 0x0F000 strncpy M_StringStartsWith M_StrCaseStr _MLIBC_ID_T_H  S_ISFIFO(m) (((m) & S_IFMT) == S_IFIFO) strstr M_ForceUppercase S_ISCHR(m) (((m) & S_IFMT) == S_IFCHR) S_IFIFO 0x01000 S_IXOTH 01 MLIBC_BLKSIZE_T_H  M_StringDuplicate S_IRUSR 0400 S_IFREG 0x08000 haystack buf_len MLIBC_TIMESPEC_H  S_IFDIR 0x04000 S_ISBLK(m) (((m) & S_IFMT) == S_IFBLK) MLIBC_INO_T_H  MLIBC_DEV_T_H  _SYS_STAT_H  m_random.c rndtable prndindex P_AddThinker EV_DoCeiling result_e P_FindSectorFromLineTag P_FindHighestCeilingSurrounding P_AddActiveCeiling P_RemoveActiveCeiling P_ActivateInStasisCeiling EV_CeilingCrushStop pastdest p_ceilng.c crushed P_RemoveThinker T_MoveCeiling T_MovePlane vld_close30ThenOpen p_doors.c P_FindLowestCeilingSurrounding vld_blazeOpen T_VerticalDoor EV_VerticalDoor vld_close vld_blazeClose EV_DoDoor vldoor_e P_SpawnDoorRaiseIn5Mins topwait vld_blazeRaise topcountdown vld_normal vld_raiseIn5Mins vld_open P_SpawnDoorCloseIn30 EV_DoLockedDoor deltax deltay A_PlayerScream A_KeenDie A_BrainPain corpsehit A_SpidRefire olddir A_Scream PIT_VileCheck braintargeton xspeed A_SkelMissile A_VileTarget actor P_SetThingPosition P_CheckMissileRange A_BabyMetal A_XScream P_TryWalk junk dirtype_t TRACEANGLE lowerFloorToLowest currentthinker DI_SOUTHEAST P_Move bangle CheckBossEnd A_FatAttack1 A_FatAttack2 A_FatAttack3 A_Chase A_Tracer NUMDIRS P_SubstNullMobj lowerAndChange P_SpawnPuff P_SetMobjState A_PainDie P_LineAttack A_BruisAttack A_TroopAttack prestep R_PointToAngle2 EV_DoFloor P_LookForPlayers raiseFloorToNearest A_BrainScream DI_SOUTHWEST raiseFloor24 exact SKULLSPEED (20*FRACUNIT) A_VileStart A_BrainAwake P_CheckSight A_VileChase A_SkelFist A_CPosAttack raiseFloor A_LoadShotgun2 newmobj soundblocks A_VileAttack P_CheckMeleeRange P_AimLineAttack DI_NORTH good A_FireCrackle DI_NORTHEAST nomissile lowerFloor A_BrainSpit DI_EAST viletryy A_BspiAttack allaround A_Fire P_LineOpening thingy vileobj turboLower numbraintargets A_Explode P_RadiusAttack A_StartFire DI_NORTHWEST seeyou raiseFloor512 A_CloseShotgun2 A_OpenShotgun2 A_PainShootSkull DI_WEST A_ReFire A_Fall raiseFloor24AndChange P_BlockThingsIterator donutRaise P_AproxDistance DI_NODIR raiseFloorCrush A_PosAttack P_UnsetThingPosition A_Hoof P_TeleportMove A_FatRaise A_Pain P_TryMove A_SargAttack P_RecursiveSound maxdist A_Look A_BrainDie A_SpawnSound A_HeadAttack A_CPosRefire A_PainAttack P_UseSpecialLine DI_SOUTH A_Metal A_CyberAttack A_BossDeath p_enemy.c A_SpawnFly A_FaceTarget A_SkullAttack P_NewChaseDir turnaround P_NoiseAlert P_DamageMobj A_SPosAttack yspeed raiseFloorTurbo FATSPREAD (ANG90/8) A_SkelWhoosh P_SpawnMissile viletryx A_BrainExplode emmiter try_ok tdir motype diags raiseToTexture opposite floorOrCeiling lastpos floortype minsize P_ChangeSector P_FindHighestFloorSurrounding getSide twoSided newspecial stair_e stairsize tsec flag p_floor.c EV_BuildStairs T_MoveFloor floor_e getSector newsecnum turbo16 P_FindNextHighestFloor floordestheight P_FindLowestFloorSurrounding build8 P_GiveBody INVULNTICS P_DropWeapon INVISTICS CF_NOCLIP hits P_GiveCard P_GiveWeapon p_inter.c P_GiveAmmo P_GiveArmor gaveammo saved __P_INTER__  CF_GODMODE thrust IRONTICS INFRATICS CF_NOMOMENTUM power card_t inflictor toucher dropped P_GivePower oldammo P_TouchSpecialThing BONUSADD 6 gaveweapon P_KillMobj P_SpawnLightFlash templine P_SpawnStrobeFlash fireflicker_t getNextSector fastOrSlow P_FindMinSurroundingLight amount T_FireFlicker bright maxtime maxlight T_StrobeFlash p_lights.c T_Glow P_SpawnFireFlicker darktime flick P_SpawnGlowingLight EV_LightTurnOn EV_StartLightStrobing T_LightFlash minlight inSync mintime brighttime EV_TurnTagLightsOff movelen secondslideline attackrange newx PTR_AimTraverse slidemo PIT_StompThing P_ThingHeightClip crunch trailx traily retry P_HitSlideLine PIT_CheckThing P_BoxOnLineSide PTR_UseTraverse thingtopslope tmdropoffz p_map.c hitcount nofit bestslideline baseaddr newy P_UseLines PIT_CheckLine P_ShootSpecialLine tmbbox leady newsubsec DEFAULT_SPECHIT_MAGIC 0x01C09C98 newlen oldside shootz deltaangle P_PathTraverse tmthing PTR_ShootTraverse onfloor tmxmove aimslope stairstep bombsource blockdist oldx oldy SpechitOverrun hitline leadx lineangle PIT_RadiusAttack usething tmflags tmymove bestslidefrac bombdamage PIT_ChangeSector isblocking P_BlockLinesIterator la_damage P_SpawnBlood secondslidefrac P_CrossSpecialLine P_SlideMove PTR_SlideTraverse crushchange thingbottomslope P_PointOnLineSide shootthing moveangle bombspot num_intercepts blockx blocky mapx mapy traverser_t PIT_AddLineIntercepts partial InterceptsMemoryOverrun earlyout ptflags xintercept PIT_AddThingIntercepts trav InterceptsOverrun yintercept maxfrac P_TraverseIntercepts p_maputl.c intercepts_overrun mapxstep bulletslope int16_array scan P_InterceptVector P_PointOnDivlineSide P_MakeDivline mapystep tmbox intercepts_overrun_t tracepositive P_RespawnSpecials P_ExplodeMissile test ptryx P_SpawnMapThing p_mobj.c FRICTION 0xe800 correct_lost_soul_bounce dummy_mobj P_CheckMissileSpawn ST_Start P_ZMovement S_StopSound P_XYMovement STOPSPEED 0x1000 P_NightmareRespawn P_SetupPsprites P_MobjThinker ptryy P_SpawnPlayerMissile T_PlatRaise p_plats.c EV_StopPlat P_RemoveActivePlat EV_DoPlat P_AddActivePlat P_ActivateInStasis P_BulletSlope A_FirePistol P_GunShot A_BFGsound A_FirePlasma A_Light1 A_Light2 A_Punch A_FireBFG A_WeaponReady WEAPONTOP 32*FRACUNIT A_FireMissile P_SetPsprite WEAPONBOTTOM 128*FRACUNIT swingy P_MovePsprites p_pspr.c DecreaseAmmo A_CheckReload P_CheckAmmo P_CalcSwing swingx accurate A_Saw swing A_FireCGun P_BringUpWeapon A_FireShotgun A_FireShotgun2 newstate ammonum LOWERSPEED FRACUNIT*6 RAISESPEED FRACUNIT*6 A_Raise A_Lower A_Light0 A_BFGSpray P_FireWeapon A_GunFlash tc_floor saveg_write_glow_t saveg_read_ceiling_t basename saveg_write_pspdef_t tc_plat saveg_write16 saveg_write_plat_t tc_door P_InitThinkers SAVEGAME_EOF 0x1d p_saveg.c saveg_read_plat_t saveg_write_think_t saveg_write_actionf_t saveg_write_floormove_t saveg_writep tc_strobe saveg_read_strobe_t saveg_read_thinker_t saveg_write_strobe_t saveg_write_player_t saveg_read_ticcmd_t padding saveg_write_ticcmd_t saveg_read_mapthing_t tc_flash saveg_read_floormove_t saveg_read_glow_t saveg_write_pad tc_ceiling tclass __mlibc_intptr specials_e saveg_write8 tc_mobj saveg_write_ceiling_t saveg_read8 saveg_readp saveg_write_mapthing_t read_vcheck saveg_read_player_t saveg_read_enum saveg_read32 saveg_read_think_t saveg_read_actionf_t tc_end tc_endspecials saveg_write_thinker_t tc_glow saveg_read_vldoor_t saveg_read_pad saveg_write_mobj_t saveg_write_vldoor_t filename_size saveg_read_pspdef_t savegamelength saveg_read_lightflash_t saveg_write_lightflash_t saveg_write_enum saveg_write32 saveg_read16 saveg_read_mobj_t P_LoadSegs ML_REJECT mapsubsector_t ML_BLOCKMAP P_InitSwitchList W_ReadLump P_LoadSideDefs R_InitSprites mapseg_t P_LoadSubsectors P_LoadLineDefs firstseg p_setup.c ML_LINEDEFS mapsidedef_t R_PrecacheLevel maplinedef_t W_GetNumForName MAX_DEATHMATCH_STARTS 10 null_sector_is_initialized mapvertex_t ML_NODES lumplen P_LoadVertexes P_LoadThings rejectpad numthings ML_SECTORS P_LoadBlockMap byte_num ML_SSECTORS totallines PadRejectArray padvalue playermask GetSectorAtNullAddress mapsector_t ML_SEGS ldef P_GroupLines ML_SIDEDEFS S_Start linebuffer P_InitPicAnims spawnthing W_ReleaseLumpNum mapnode_t minlength null_sector Z_FreeTags ML_LABEL P_LoadSectors P_LoadNodes ML_THINGS ML_VERTEXES P_LoadReject P_SpawnSpecials W_LumpLength bytenum P_CrossSubsector P_DivlineSide sightcounts divl sightzstart p_sight.c bitnum bspnum P_InterceptVector2 P_CrossBSPNode strace basepic DONUT_FLOORHEIGHT_DEFAULT 0x00000000 R_CheckTextureNumForName EV_DoDonut startname p_spec.c istexture anim_t tmp_s3_floorpic P_UpdateSpecials EV_Teleport first numpics DONUT_FLOORPIC_DEFAULT 0x16 pillar_sector heightlist animdefs linespeciallist tmp_s3_floorheight endname P_PlayerInSpecialSector P_ChangeSwitchTexture MAXANIMS 32 numlinespecials MAX_ADJOINING_SECTORS 20 currentheight linenum lastanim DonutOverrun currentSector MAXLINEANIMS 64 numflats animdef_t texBot texMid P_StartButton switchlist_t numswitches name1 name2 useAgain switchlist p_switch.c alphSwitchList texTop p_telept.c oldz P_PlayerThink P_AllocateThinker P_RunThinkers p_tick.c P_MovePlayer ANG5 (ANG90/18) newweapon onground MAXBOB 0x100000 P_DeathThink P_CalcHeight P_Thrust INVERSECOLORMAP 32 p_user.c R_FindPlane tspan R_StoreWallRange angle2 R_PointToAngle clippass R_ClipPassWallSegment bspcoord clipsolid R_ClipSolidWallSegment R_AddLine newend MAXSEGS 32 R_PointOnSide R_Subsector R_ClearDrawSegs R_ClearClipSegs R_CheckBBox cliprange_t boxpos checkcoord R_AddSprites solidsegs R_RenderBSPNode r_bsp.c boxx boxy Z_ChangeTag2 firstpatch texturecompositesize maxoff mpatch patchcount R_InitSpriteLumps obsolete originy R_DrawColumnInCache spritepresent texturepresent masked numtextures1 numtextures2 originx flatmemory cacheheight GenerateTextureHashTable texturecolumnofs textures_hashtable R_InitTextures R_GetColumn patchlookup R_InitData collump texpatch_t mappatch_t r_data.c numtextures texturecomposite nummappatches lastpatch colofs texturewidthmask lastflat spritememory R_GenerateLookup R_InitFlats realpatch texturememory stepdir R_InitColormaps maxoff2 temp1 temp2 temp3 totalwidth name_p maptex texture_s patchcol maptex1 texnum namet texturecolumnlump W_LumpNameHash R_GenerateComposite numpatches flatpresent maptexture_t directory maptex2 fracstep V_UseBuffer SBARHEIGHT 32 R_DrawTranslatedColumnLow R_DrawColumnLow R_DrawSpan R_InitBuffer FUZZOFF (SCREENWIDTH) R_DrawSpanLow FUZZTABLE 50 viewimage R_DrawColumn background_buffer fuzzpos MAXHEIGHT 832 R_DrawTranslatedColumn dscount xtemp ylookup dccount R_DrawFuzzColumn MAXWIDTH 1120 ytemp r_draw.c translations fuzzoffset R_DrawFuzzColumnLow R_InitTranslationTables walllights R_ScaleFromGlobalAngle R_ClearPlanes angleb R_InitTables R_InitLightTables anglea R_InitPointToAngle R_SetupFrame sineb focallength framecount R_ClearSprites sinea R_InitPlanes FIELDOFVIEW 2048 SlopeDiv r_main.c R_PointOnSegSide DISTMAP 2 cosadj R_PointToDist R_AddPointToBox nodenum visangle R_DrawPlanes R_InitSkyMap setdetail R_DrawMasked R_InitTextureMapping setblocks R_MakeSpans cacheddistance spanstop baseyscale R_CheckPlane unionh unionl visplanes planeheight openings ceilingfunc basexscale intrh spanstart MAXVISPLANES 128 MAXOPENINGS SCREENWIDTH*64 cachedxstep planezlight lastvisplane intrl R_MapPlane cachedystep cachedheight r_plane.c offsetangle R_DrawMaskedColumn r_segs.c rw_midtexturemid HEIGHTBITS 12 bottomfrac rw_bottomtexturemid pixhighstep rw_scale topfrac distangle texturecolumn worldbottom worldhigh lightnum bottomstep rw_centerangle worldtop vtop HEIGHTUNIT (1<<HEIGHTBITS) sineval R_RenderMaskedSegRange maskedtexture worldlow pixlowstep R_RenderSegLoop rw_offset pixhigh pixlow rw_toptexturemid rw_scalestep topstep r_sky.c newvissprite tr_y flipped R_DrawPlayerSprites rotation avis basetexturemid R_InstallSpriteLump sprtemp lowscale clipbot namelist unsorted R_DrawVisSprite r_things.c R_DrawPSprite patched spritelights bottomscreen R_SortVisSprites R_InitSpriteDefs R_DrawSprite bestscale BASEYCENTER 100 R_NewVisSprite spritename R_ProjectSprite MINZ (FRACUNIT*4) cliptop overflowsprite tr_x maxframe sha1_context_s K4 0xCA62C1D6L X(a) do { *p++ = hd->h ##a >> 24; *p++ = hd->h ##a >> 16; *p++ = hd->h ##a >> 8; *p++ = hd->h ##a; } while(0) rol(x,n) ( ((x) << (n)) | ((x) >> (32-(n))) ) SHA1_UpdateInt32 SHA1_Update digest sha1_context_t K1 0x5A827999L K3 0x8F1BBCDCL SHA1_UpdateString K2 0x6ED9EBA1L assert(assertion) ((void)((assertion) || (__assert_fail(#assertion, __FILE__, __LINE__, __func__), 0))) R(a,b,c,d,e,f,k,m) do { e += rol( a, 5 ) + f( b, c, d ) + k + m; b = rol( b, 30 ); } while(0) sha1.c inbuf assert Transform F3(x,y,z) ( ( x & y ) | ( z & ( x | y ) ) ) F2(x,y,z) ( x ^ y ^ z ) SHA1_Init F1(x,y,z) ( z ^ ( x & ( y ^ z ) ) ) F4(x,y,z) ( x ^ y ^ z ) SHA1_Final M(i) ( tm = x[i&0x0f] ^ x[(i-14)&0x0f] ^ x[(i-8)&0x0f] ^ x[(i-3)&0x0f] , (x[i&0x0f] = rol(tm,1)) ) _ASSERT_H  inlen SOUND(name,priority) { NULL, name, priority, NULL, -1, -1, 0, 0, -1, NULL } sounds.c MUSIC(name) { name, 0, NULL, NULL } SOUND_LINK(name,priority,link_id,pitch,volume) { NULL, name, priority, &S_sfx[link_id], pitch, volume, 0, 0, -1, NULL } doom1_par_times num_captured_stats statdump.c StatDump doom2_par_times MAX_CAPTURES 32 st_multicon_t STlib_initPercent STlib_initBinIcon STlib_init V_CopyRect oldinum st_lib.c STlib_initNum STlib_initMultIcon sttminus __STLIB__  STlib_updateMultIcon oldnum STlib_updateBinIcon STlib_updateNum STlib_updatePercent numdigits STlib_drawNum st_binicon_t st_number_t st_percent_t oldval ST_doRefresh ST_TURNCOUNT (1*TICRATE) ST_AMMO0Y 173 ST_FRAGSWIDTH 2 st_oldhealth ST_initData ST_MAXAMMO0HEIGHT 5 ST_MAPTITLEY 0 ST_AMMOY 171 st_firsttime ST_WEAPON4Y 181 st_randomnumber st_chatstateenum_t ST_GODFACE (ST_NUMPAINFACES*ST_FACESTRIDE) ST_KEY0HEIGHT 5 w_frags ST_AMMO1X 288 ST_WEAPON2Y 172 ST_DETHX 109 w_faces ST_MAPTITLEX (SCREENWIDTH - ST_MAPWIDTH * ST_CHATFONTWIDTH) st_msgcounter STARTBONUSPALS 9 ST_EVILGRINOFFSET (ST_OUCHOFFSET + 1) ST_RAMPAGEOFFSET (ST_EVILGRINOFFSET + 1) ST_MAXAMMO3X 314 ST_MSGTEXTX 0 ST_DEADFACE (ST_GODFACE+1) largeammo st_facecount ST_AMMO3X 288 w_arms ST_KEY2X 239 ST_AMMO1WIDTH ST_AMMO0WIDTH ST_FRAGSY 171 lastattackdown ST_MSGHEIGHT 1 ST_MSGWIDTH 52 ST_OUTTEXTX 0 ST_calcPainOffset ST_NUMEXTRAFACES 2 ST_ARMSBGX 104 musnum ST_KEY0Y 171 w_maxammo lastcalc ST_MAXAMMO3Y 185 ST_updateFaceWidget StartChatState ST_drawWidgets st_palette diffang w_health ST_unloadGraphics ST_X2 104 ST_AMMO2Y 191 ST_NUMTURNFACES 2 ST_KEY0WIDTH 8 ST_AMMOWIDTH 3 RADIATIONPAL 13 ST_unloadData ST_MAXAMMO0Y 173 NUMREDPALS 8 GetChatState ST_DETHY 191 ST_FX 143 ST_STRAIGHTFACECOUNT (TICRATE/2) FirstPersonState ST_MAXAMMO1Y 179 ST_KEY2WIDTH ST_KEY0WIDTH ST_WEAPON5Y 181 ST_WEAPON5X 134 ST_AMMO2X 288 ST_MUCHPAIN 20 w_ammo st_statusbaron ST_ARMORWIDTH 3 shortnum ST_ARMSBGY 168 ST_NUMPAINFACES 5 ST_FACESTRIDE (ST_NUMSTRAIGHTFACES+ST_NUMTURNFACES+ST_NUMSPECIALFACES) ST_MAXAMMO3WIDTH ST_MAXAMMO0WIDTH w_armsbg ST_ARMSX 111 ST_loadCallback ST_FY 169 ST_loadGraphics faceback ST_MAXAMMO2WIDTH ST_MAXAMMO0WIDTH NUMBONUSPALS 4 ST_ARMSYSPACE 10 st_fragscount ST_TOGGLECHAT KEY_ENTER ST_WEAPON4X 122 ST_MAXAMMO0X 314 ST_MAXAMMO1X 314 ST_diffDraw ST_KEY1Y 181 w_ready st_fragson st_armson ST_WEAPON1X 122 st_notdeathmatch ST_WEAPON3X 110 ST_KEY0X 239 AutomapState ST_ARMSXSPACE 12 st_oldchat ST_AMMO3Y 185 lu_palette ST_FACEPROBABILITY 96 ST_loadUnloadGraphics ST_WEAPON2X 134 ST_AMMO0HEIGHT 6 ST_HEALTHX 90 ST_ARMORX 221 ST_OUTTEXTY 6 ST_AMMOX 44 ST_ARMSY 172 ST_AMMO1Y 179 ST_AMMO0WIDTH 3 ST_OUTWIDTH 52 ST_NUMFACES (ST_FACESTRIDE*ST_NUMPAINFACES+ST_NUMEXTRAFACES) ST_MSGTEXTY 0 st_cursoron ST_OUCHOFFSET (ST_TURNOFFSET + ST_NUMTURNFACES) ST_doPaletteStuff ST_unloadCallback st_clock ST_KEY1WIDTH ST_KEY0WIDTH ST_RAMPAGEDELAY (2*TICRATE) st_stateenum_t ST_HEALTHWIDTH 3 ST_MAPHEIGHT 1 tallpercent ST_WEAPON1Y 172 ST_refreshBackground doevilgrin badguyangle ST_AMMO0X 288 ST_FACESX 143 ST_OUTHEIGHT 1 st_stuff.c w_keyboxes ST_KEY1X 239 ST_WPNSX 109 tallnum ST_HEALTHY 171 ST_MAXAMMO2X 314 ST_updateWidgets ST_WEAPON3Y 181 ST_loadData st_gamestate ST_Stop ST_OUCHCOUNT (1*TICRATE) ST_NUMSPECIALFACES 3 st_chatstate ST_AMMO2WIDTH ST_AMMO0WIDTH ST_KEY2Y 191 ST_X 0 ST_NUMSTRAIGHTFACES 3 st_chat ST_createWidgets STARTREDPALS 1 oldweaponsowned ST_MAXAMMO2Y 191 w_armor ST_FACESY 168 ST_TURNOFFSET (ST_NUMSTRAIGHTFACES) ST_MAXAMMO0WIDTH 3 st_faceindex ST_MAXAMMO1WIDTH ST_MAXAMMO0WIDTH ST_FRAGSX 138 facenum load_callback_t st_stopped ST_EVILGRINCOUNT (2*TICRATE) ST_WEAPON0X 110 ST_AMMO3WIDTH ST_AMMO0WIDTH WaitDestState ST_WEAPON0Y 172 ST_WPNSY 191 ST_ARMORY 171 ST_TALLNUMWIDTH (tallnum[0]->width) snd_SfxVolume S_AdjustSoundParams listener sfx_id s_sound.c S_StopChannel S_ATTENUATOR ((S_CLIPPING_DIST - S_CLOSE_DIST) >> FRACBITS) mus_playing m_id S_StopMusic spmus NORM_SEP 128 S_CLOSE_DIST (200 * FRACUNIT) audible S_GetChannel NORM_PITCH 128 mus_paused musicnum approx_dist mnum channel_t origin_p S_CLIPPING_DIST (1200 * FRACUNIT) NORM_PRIORITY 64 S_MusicPlaying origin S_Shutdown S_STEREO_SWING (96 * FRACUNIT) tables.c patchclip_callback bits_per_pixel V_DrawShadowedPatch palette_type destx desty MOUSE_SPEED_BOX_HEIGHT 9 I_GetPaletteIndex xmax V_DrawTLPatch V_DrawRawScreen V_LoadXlaTable redline_x V_DrawVertLine desttop2 V_DrawBox lbmname V_DrawFilledBox vres WritePCXfile encoding V_DrawAltTLPatch V_DrawHorizLine manufacturer format ymax usemouse bordercolor xmin buf1 vpatchclipfunc_t pcx_t color_planes filler xlatab dest_screen v_video.c white bgcolor V_SetPatchClipCallback srcx srcy black yellow linelen MOUSE_SPEED_BOX_WIDTH 120 V_LoadTintTable V_DrawXlaPatch bytes_per_line reserved hres box_x box_y ymin original_speed WI_initVariables WI_initNoState WI_initShowNextLoc SP_FRAGS 6 stillticking WI_slamBackground sp_secret WI_drawNetgameStats fontwidth cnt_par killers WI_drawAnimatedBack ANIM_RANDOM SP_TIMEY (SCREENHEIGHT-32) WI_drawNum WI_updateNoState WI_initDeathmatchStats WI_initStats WI_updateDeathmatchStats victims sucks SP_TIME 8 WI_drawShowNextLoc WI_initNetgameStats SP_PAR ST_TIME dm_state WI_drawTime animenum_t SP_SECRET 4 DM_TOTALSX 269 WI_unloadCallback DM_SPACINGX 40 WI_loadCallback NG_STATSX (32 + SHORT(star->width)/2 + 32*!dofrags) finished ANIM(type,period,nanims,x,y,nexttic) { (type), (period), (nanims), { (x), (y) }, (nexttic), 0, { NULL, NULL, NULL }, 0, 0, 0, 0 } dm_frags splat WI_fragSum SP_STATSY 50 cnt_pause epsd2animinfo WI_drawOnLnode StatCount entering DM_VICTIMSY 50 fsum epsd1animinfo cnt_time lastdrawn fits NG_STATSY 50 ng_state NUMMAPS 9 SP_TIMEX 16 NG_SPACINGX 64 DM_VICTIMSX 5 firstrefresh SP_STATSX 50 sp_state NUMEPISODES 4 period WI_drawPercent SP_KILLS 0 WI_initAnimatedBack lnames WI_checkForAccelerate bstar DM_KILLERSY 100 colon WI_Responder DM_KILLERSX 10 dofrags NUMANIMS WI_unloadData WI_updateNetgameStats wiminus WI_updateShowNextLoc dm_totals WI_drawEL WI_drawDeathmatchStats WI_drawNoState SP_PAUSE 1 timepatch acceleratestage WI_drawStats WI_TITLEY 2 WI_drawLF DM_MATRIXY 68 epsd0animinfo WI_SPACINGY 33 cnt_frags SHOWNEXTLOCDELAY 4 ANIM_ALWAYS lnodes WI_updateAnimatedBack cnt_kills ANIM_LEVEL WI_loadData nanims DM_MATRIXX 42 wbstartstruct plrs bcnt WI_loadUnloadData NUMCMAPS wi_stuff.c snl_pointeron cnt_items WI_updateStats SP_ITEMS 2 cnt_secret realloc sha1_context ChecksumAddLump num_open_wadfiles w_checksum.c GetFileNumber wad_file_classes w_file.c W_CloseFile W_OpenFile stdc_wad_file buffer_len W_Read w_main.c W_NWT_MERGE_FLATS 0x2 W_MERGE_H  W_NWT_MERGE_SPRITES 0x1 header fileinfo I_EndRead newnumlumps filelump_t I_BeginRead identification filerover lumphash w_wad.c unique_lumps startlump wadinfo_t newlumpinfo calloc ExtendLumpInfo filepos W_NumLumps lump_p infotableofs nextlumpnum Z_ChangeUser mainzone Z_ClearZone user Z_ZoneSize lowtag Z_FreeMemory z_zone.c newblock Z_FileDumpHeap hightag blocklist memzone_t Z_DumpHeap memblock_s memblock_t ZONEID 0x1d4a11 MEM_ALIGN sizeof(void *) MINFRAGMENT 64 W_StdC_CloseFile stdc_wad_file_t W_StdC_Read stdc_wad w_file_stdc.c W_StdC_OpenFile __MLIBC_O_DSYNC 0x0800 O_NDELAY __MLIBC_O_NONBLOCK _ABIBITS_ABI_H  __MLIBC_O_RDWR 3 F_SETLK 8 __MLIBC_O_NONBLOCK 0x0400 AT_FDCWD -100 O_EXEC __MLIBC_O_EXEC O_NOCTTY __MLIBC_O_NOCTTY at_to_doom O_APPEND __MLIBC_O_APPEND F_GETLK 7 O_NOFOLLOW __MLIBC_O_NOFOLLOW _ABIBITS_FCNTL_H  O_EXCL __MLIBC_O_EXCL O_DIRECTORY __MLIBC_O_DIRECTORY F_SETFL 6 __MLIBC_O_TRUNC 0x0200 __MLIBC_O_WRONLY 5 AT_EMPTY_PATH 1 __MLIBC_O_DIRECTORY 0x0020 F_SETOWN 11 O_WRONLY __MLIBC_O_WRONLY F_GETFL 5 POSIX_FADV_NORMAL 1 __MLIBC_O_SEARCH 4 F_SETLKW 9 shiftdown O_CREAT __MLIBC_O_CREAT F_UNLCK 2 F_WRLCK 3 DG_GetKey pressed O_TRUNC __MLIBC_O_TRUNC shiftxform __MLIBC_O_EXEC 1 GetTypedChar POSIX_FADV_WILLNEED 5 __MLIBC_O_ACCMODE 0x0007 __MLIBC_O_NOFOLLOW 0x0100 O_ACCMODE __MLIBC_O_ACCMODE UpdateShiftStatus __MLIBC_O_CLOEXEC 0x4000 F_GETOWN 10 F_SETFD 4 F_DUPFD 1 FD_CLOEXEC 1 POSIX_FADV_DONTNEED 4 POSIX_FADV_SEQUENTIAL 2 F_GETFD 3 POSIX_FADV_RANDOM 6 __MLIBC_O_RDONLY 2 __MLIBC_O_APPEND 0x0008 POSIX_FADV_NOREUSE 3 O_DSYNC __MLIBC_O_DSYNC AT_SYMLINK_NOFOLLOW 4 F_RDLCK 1 __I_SCALE__  I_InitInput i_input.c __MLIBC_O_EXCL 0x0040 O_CLOEXEC __MLIBC_O_CLOEXEC O_RDWR __MLIBC_O_RDWR __MLIBC_O_CREAT 0x0010 __MLIBC_O_NOCTTY 0x0080 O_SEARCH __MLIBC_O_SEARCH AT_SYMLINK_FOLLOW 2 AT_EACCESS 512 O_NONBLOCK __MLIBC_O_NONBLOCK F_DUPFD_CLOEXEC 2 TranslateKey __MLIBC_O_SYNC 0x2000 O_SYNC __MLIBC_O_SYNC I_GetEvent O_RDONLY __MLIBC_O_RDONLY AT_REMOVEDIR 8 O_RSYNC __MLIBC_O_RSYNC __MLIBC_O_RSYNC 0x1000 dots_on x_offset_end grabmouse_callback_t transp rcsid GFX_RGB565_R(color) ((0xF800 & color) >> 11) x_offset cmap_to_rgb565 $Id: i_x.c,v 1.6 1997/02/03 22:45:10 b1 Exp $ __mlibc_uint16 GFX_RGB565(r,g,b) ((((r & 0xF8) >> 3) << 11) | (((g & 0xFC) >> 2) << 5) | ((b & 0xF8) >> 3)) xres bool _Bool in_pixels line_in I_ShutdownGraphics DG_DrawFrame blue line_out GFX_RGB565_B(color) (0x001F & color) xres_virtual GFX_RGB565_G(color) ((0x07E0 & color) >> 5) _STDBOOL_H  DG_SetWindowTitle cmap_to_fb I_VideoBuffer_FB true 1 rgb565_palette uint16_t col_t y_offset FB_ScreenInfo FB_BitField yres false 0 green yres_virtual __bool_true_false_are_defined 1 s_Fb fb_scaling i_video.c DG_Init doomgeneric.c _GLIBCXX_GTHREAD_USE_WEAK 0 __cpp_aggregate_nsdmi 201304 _ZSt3absd _ZSt3absg _GLIBCXX_HAVE_ENOTRECOVERABLE 1 _ZSt3absl _GLIBCXX_INCLUDE_NEXT_C_HEADERS _ZSt3absn _ZSt3absx _GLIBCXX_HAVE_ACOSL 1 _GLIBCXX_HAVE_SINHL 1 _GLIBCXX_DEPRECATED __attribute__ ((__deprecated__)) _GLIBCXX_USE_C99_MATH _GLIBCXX11_USE_C99_MATH _GLIBCXX_HAVE_STRINGS_H 1 WINDOW_FLAGS_SNAP_TO_BOTTOM 0x2 _GLIBCXX_PSEUDO_VISIBILITY(V)  SYS_STAT 18 _GLIBCXX11_USE_C99_STDLIB 1 __DBL_EPSILON__ double(2.22044604925031308084726333618164062e-16L) _GLIBCXX_USE_C99_STDIO _GLIBCXX11_USE_C99_STDIO KEY_ARROW_DOWN 269 _GLIBCXX_TXN_SAFE  _GLIBCXX_HAVE_EPROTO 1 _GLIBCXX_HAVE_FLOORF 1 SYS_OPEN 5 _GLIBCXX_HAVE_COSL 1 _GLIBCXX_HAVE_LIMIT_FSIZE 1 __cpp_alias_templates 200704 _GLIBCXX_HAVE_DLFCN_H 1 NULL __null WINDOW_EVENT_MOUSEUP 3 strtoll KEY_F1 256 _GLIBCXX_USE_C99_COMPLEX _GLIBCXX11_USE_C99_COMPLEX __MLIBC_STATIC_ASSERT(c,text) static_assert(c, text) __DBL_DENORM_MIN__ double(4.94065645841246544176568792868221372e-324L) _GLIBCXX_HAVE_COSHF 1 _GLIBCXX_HAVE_HYPOTF 1 _GLIBCXX_VERBOSE 1 WindowPaintHandler _GLIBCXX_HAVE_MBSTATE_T 1 senderPID _BSD_PTRDIFF_T_  _GLIBCXX_HAVE_EOVERFLOW 1 UpdateWindow _GLIBCXX_HAVE_ECANCELED 1 atoll KEY_STATE_CONTROL 8 _GLIBCXX_HAVE_TGMATH_H 1 lastPressedWidget KEY_ARROW_UP 266 SYS_MAP_FB 14 __STDC_LIMIT_MACROS _GLIBCXX_HAVE_POWF 1 SYS_READ 3 SYS_RENDER_WINDOW 27 DESKTOP_EVENT 0xBEEF KEY_F5 260 _GLIBCXX_SYNCHRONIZATION_HAPPENS_BEFORE(A)  IPC_H  atol SYSCALL_H  _GLIBCXX_HAVE_WCHAR_H 1 _GLIBCXX_HAVE_FENV_H 1 doomgeneric_lemon.cpp recieverPID _GLIBCXX_HAVE_QUICK_EXIT 1 getenv __cpp_variable_templates 201304 _GLIBCXX_BITS_STD_ABS_H  KEY_CONTROL 272 _GLIBCXX17_DEPRECATED  __cpp_hex_float 201603 KEY_STATE_SHIFT 2 _GLIBCXX_NOEXCEPT_QUAL  wctomb _GLIBCXX_END_NAMESPACE_VERSION  primaryBuffer _GLIBCXX_USE_C99_WCHAR _GLIBCXX11_USE_C99_WCHAR _GLIBCXX_HAVE_ETIMEDOUT 1 tolower s_KeyQueueWriteIndex SYS_CREATE 8 ReceiveMessage KEY_F6 261 _GLIBCXX_LONG_DOUBLE_COMPAT _GLIBCXX_NOEXCEPT noexcept _GLIBCXX_DEFAULT_ABI_TAG _GLIBCXX_ABI_TAG_CXX11 _GLIBCXX_HAVE_VFWSCANF 1 _GLIBCXX_BEGIN_NAMESPACE_ALGO  _GLIBCXX_HAVE_ATANF 1 __cpp_lambdas 200907 _GLOBAL__sub_I_window _GLIBCXX_CONST __attribute__ ((__const__)) _GLIBCXX_HAVE_ENOTSUP 1 _GLIBCXX_HAVE_SYS_STATVFS_H 1 _ZN4ListIP6WidgetED4Ev _GLIBCXX_NORETURN __attribute__ ((__noreturn__)) s_KeyQueue _GLIBCXX_BEGIN_NAMESPACE_LDBL_OR_CXX11 _GLIBCXX_BEGIN_NAMESPACE_CXX11 _GLIBCXX_HOSTED 1 strtoull SYS_EXEC 2 SURFACE_H  _GLIBCXX_CSTDLIB 1 _GLIBCXX11_USE_C99_STDIO 1 __cpp_constexpr 201304 SYS_WAIT_PID 38 _GLIBCXX14_CONSTEXPR constexpr __cpp_generic_lambdas 201304 _GLIBCXX_HAVE_ETXTBSY 1 __cpp_digit_separators 201309 SwapWindowBuffers KEY_SHIFT 270 ownerPID remove_at _GLIBCXX_HAVE_STRTOLD 1 _GLIBCXX_PACKAGE_TARNAME "libstdc++" SYS_CLOSE 6 linePadding 7lldiv_t _GLIBCXX_END_EXTERN_C } KEY_ARROW_RIGHT 268 _GLIBCXX_USE_FLOAT128 1 _GLIBCXX_HAVE_MODFF 1 __GLIBCXX_TYPE_INT_N_0 __int128 KEY_BACKSPACE '\b' add_front _Z17SwapWindowBuffersP6Window __N(msgid) (msgid) _GLIBCXX_HAVE_SYS_TIME_H 1 SYS_GET_VIDEO_MODE 31 _GLIBCXX_HAVE_LOCALE_H 1 __cpp_variadic_templates 200704 WINDOW_FLAGS_MINIMIZED 0x4 _ZN9__gnu_cxx3divExx WINDOW_EVENT_KEY 1 _GLIBCXX_TXN_SAFE_DYN  _GLIBCXX_HAVE_LIMIT_AS 1 SYS_READDIR 33 SYS_UPTIME 30 _GLIBCXX11_USE_C99_MATH 1 _GLIBCXX_PURE __attribute__ ((__pure__)) _GLIBCXX_NAMESPACE_LDBL_OR_CXX11 _GLIBCXX_NAMESPACE_CXX11 _GLIBCXX_HAVE_EWOULDBLOCK 1 llabs WINDOW_EVENT_MOUSEMOVE 6 5div_t _GLIBCXX_STDIO_SEEK_CUR 1 vector2i_t __cpp_range_based_for 200907 decltype(nullptr) _GLIBCXX_HAVE_HYPOT 1 strcpy mblen handle_t __static_initialization_and_destruction_0 KEY_ENTER '\n' _GLIBCXX_PACKAGE_NAME "package-unused" SYS_UNAME 32 _ZN4ListIP6WidgetE8get_backEv _GLIBCXX_HAVE_DIRENT_H 1 _GLIBCXX_STDIO_EOF -1 _GLIBCXX_BEGIN_NAMESPACE_LDBL  _GLIBCXX_ABI_TAG_CXX11 __attribute ((__abi_tag__ ("cxx11"))) __STDC_CONSTANT_MACROS _GLIBCXX_HAVE_LOGF 1 _GLIBCXX_FAST_MATH 0 __cpp_sized_deallocation 201309 _GLIBCXX_HAVE_SQRTF 1 _KEY_ESCAPE 27 _GLIBCXX_HAVE_HYPOTL 1 _GLIBCXX_END_NAMESPACE_LDBL_OR_CXX11 _GLIBCXX_END_NAMESPACE_CXX11 _GLIBCXX_HAVE_VWSCANF 1 __cpp_decltype 200707 _GLIBCXX_HAVE_SYS_IOCTL_H 1 _GLIBCXX_HAVE_MODFL 1 SYS_DESKTOP_GET_WINDOW_COUNT 25 _GLIBCXX98_USE_C99_STDLIB 1 _GLIBCXX_HAVE_LIMIT_DATA 1 seconds __cpp_ref_qualifiers 200710 _GLIBCXX_HAVE_FMODL 1 _GLIBCXX_HAVE_STDINT_H 1 clear keyCode strtoul _GLIBCXX_CONSTEXPR constexpr _GLIBCXX_HAVE_SINCOS 1 _GLIBCXX_NAMESPACE_LDBL  SYS_NANO_SLEEP 39 RGBAColour _ZN10win_info_tC2Ev _GLIBCXX_HAVE_AS_SYMVER_DIRECTIVE 1 syscall(call,arg0,arg1,arg2,arg3,arg4) asm volatile("int $0x69" :: "a"(call), "b"(arg0), "c"(arg1), "d"(arg2), "S"(arg3), "D"(arg4)) SYS_SLEEP 7 _GLIBCXX_HAVE_WCTYPE_H 1 SYS_CHMOD 16 _ZSt3abse _ZN4ListIP6WidgetE9get_frontEv _GLIBCXX_HAVE_EXPF 1 _GLIBCXX_EXTERN_TEMPLATE 1 __priority _GLIBCXX_OS_DEFINES 1 _GLIBCXX_HAVE_STDBOOL_H 1 _GLIBCXX_HAVE_LDEXPF 1 __cpp_raw_strings 200710 add_back _GLIBCXX_USE_INT128 1 _GLIBCXX_THROW(_EXC)  _GLIBCXX_HAVE_POWL 1 _Z13DestroyWindowP6Window __cpp_nsdmi 200809 LT_OBJDIR ".libs/" operator[] __cpp_static_assert 200410 _Exit strtof _GLIBCXX_HAVE_TANHL 1 _GLIBCXX_USE_DEPRECATED 1 SYS_DESKTOP_GET_WINDOW 24 replace_at _Z12UpdateWindowP6Window offsetof(TYPE,MEMBER) __builtin_offsetof (TYPE, MEMBER) wcstombs __DBL_MAX__ double(1.79769313486231570814527423731704357e+308L) _ZN4ListIP6WidgetE8add_backES1_ _GLIBCXX_HAVE_MODF 1 __float128 __cpp_attributes 200809 KEY_F4 259 SYS_GET_CWD 37 _GLIBCXX_HAVE_LOG10F 1 _GLIBCXX_X86_RDRAND 1 _T_PTRDIFF_  _GXX_NULLPTR_T  __cplusplus 201402L _GLIBCXX_HAVE_UTIME_H 1 _GLIBCXX_CXX_CONFIG_H 1 _GLIBCXX_HAVE_INTTYPES_H 1 _GLIBCXX_BEGIN_NAMESPACE_CONTAINER  SYS_PWRITE 41 __mlibc_uint64 __need_ptrdiff_t __initialize_p _GLIBCXX_HAVE_ASINF 1 surface SYS_CREATE_DESKTOP 17 _GLIBCXX_HAVE_LOG10L 1 KEY_F2 257 OnPaint secondaryBuffer _ZN4ListIP6WidgetE9remove_atEj _GLIBCXX_USE_C99_INTTYPES_TR1 1 SYS_MMAP 35 s_KeyQueueReadIndex _GLIBCXX_HAVE_SYS_TYPES_H 1 _GLIBCXX_USE_C99_STDINT_TR1 1 _GLIBCXX_HAVE_SINCOSF 1 __cpp_threadsafe_static_init 200806 _GLIBCXX_HAVE_LC_MESSAGES 1 _GLIBCXX_NAMESPACE_CXX11 __cxx11:: _GLIBCXX_HAVE_COSHL 1 _GLIBCXX_STD_C std SYS_PREAD 40 SYS_LSEEK 19 mbtowc _GLIBCXX_USE_C99 1 depth _GLIBCXX_HAVE_TANHF 1 _GLIBCXX_HAVE_ENDIAN_H 1 _GLIBCXX_HAVE_VSWSCANF 1 __cpp_delegating_constructors 200604 __GXX_EXPERIMENTAL_CXX0X__ 1 _GLIBCXX_USE_WCHAR_T 1 _GLIBCXX98_USE_C99_STDIO 1 SYS_SET_FS_BASE 34 rgba_colour_t _ANSI_STDDEF_H  _GLIBCXX_THROW_OR_ABORT(_EXC) (throw (_EXC)) _GLIBCXX_HAVE_LOGL 1 keyData _GLIBCXX_HAVE_AT_QUICK_EXIT 1 _GLIBCXX17_CONSTEXPR  _GLIBCXX_USE_DUAL_ABI 1 qsort _GLIBCXX_PACKAGE_URL "" _GLIBCXX_INLINE_VERSION 0 __cpp_initializer_lists 200806 _GLIBCXX_BEGIN_NAMESPACE_VERSION  _GLIBCXX_HAVE_ATAN2F 1 _T_PTRDIFF  _ZN4ListIP6WidgetEixEj addKeyToQueue 6ldiv_t _GLIBCXX_NOTHROW _GLIBCXX_USE_NOEXCEPT __cpp_rvalue_reference 200610 __GLIBCXX_BITSIZE_INT_N_0 128 _GLIBCXX_HAVE_ECHILD 1 WINDOW_EVENT_CLOSE 5 _PTRDIFF_T_DECLARED  _GLIBCXX_HAVE_INT64_T 1 _GLIBCXX_HAVE_ASINL 1 ListNode<Widget*> KEY_F3 258 _GLIBCXX_HAVE_ATANL 1 KEY_ALT 271 _GLIBCXX_HAVE_COSF 1 _GLIBCXX_HAVE_SYS_PARAM_H 1 __GXX_RTTI 1 _GLIBCXX_SYNCHRONIZATION_HAPPENS_AFTER(A)  DESKTOP_EVENT_KEY 0x1BEEF __cpp_inheriting_constructors 201511 __gnu_cxx _GLIBCXX_HAVE_ENODATA 1 _GLIBCXX_HAVE_TANF 1 bool _GCC_PTRDIFF_T  _GLIBCXX_STDIO_SEEK_END 2 _GLIBCXX_HAVE_STRTOF 1 _GLIBCXX_USE_CXX11_ABI 1 long double _GLIBCXX_HAVE_FMODF 1 _GLIBCXX_HAVE_FREXPL 1 SYS_GRANT_PTY 36 memcpy_optimized SYS_WRITE 4 windowInfo _GLIBCXX_CPU_DEFINES 1 get_front __STDC_CONSTANT_MACROS  _ZN4ListIP6WidgetE6get_atEj __cpp_decltype_auto 201304 _GLIBCXX_HAVE_ATTRIBUTE_VISIBILITY 1 _GLIBCXX17_INLINE  bsearch _GLIBCXX_FULLY_DYNAMIC_STRING 0 _GLIBCXX_HAVE_LDEXPL 1 _GLIBCXX_HAVE_SINHF 1 __cpp_rtti 199711 long long unsigned int _ZN4ListIP6WidgetEC4Ev surface_t __PTRDIFF_T  _GTHREAD_USE_MUTEX_TIMEDLOCK 1 _GLIBCXX_USE_ALLOCATOR_NEW 1 KEY_F9 264 _GLIBCXX_NOEXCEPT_PARM  KEY_STATE_ALT 4 _ZSt3absf SYS_CHDIR 12 doomKey _GLIBCXX_STDLIB_H 1 _GLIBCXX_HAVE_SYS_RESOURCE_H 1 __DEPRECATED 1 WINDOW_EVENT_MOUSEDOWN 2 __cpp_user_defined_literals 200809 FB_H  mousePos DESKTOP_EVENT_KEY_RELEASED 0x2BEEF _GLIBCXX_PACKAGE_STRING "package-unused version-unused" _GLIBCXX_HAVE_ENOLINK 1 _GLIBCXX_USE_CONSTEXPR constexpr __cxx11 _ZSt3divll quot KEY_ARROW_LEFT 267 ___int_ptrdiff_t_h  SYS_MOUNT 21 _GLIBCXX_END_NAMESPACE_LDBL  ~List _GLIBCXX_HAVE_STDALIGN_H 1 _GLIBCXX_HAVE_SYS_UIO_H 1 __cpp_exceptions 199711 _GLIBCXX_HAVE_SLEEP 1 SYS_ALLOC 15 _Z14ReceiveMessageP13ipc_message_t _GLIBCXX_WEAK_DEFINITION  __cpp_unicode_literals 200710 _GLIBCXX_HAVE_TANL 1 get_back _GLIBCXX_HAVE_FABSL 1 KEY_TAB '\t' _GLIBCXX_HAVE_ATAN2L 1 _GLIBCXX_HAVE_SINF 1 get_at SYS_GETPID 20 _GCC_MAX_ALIGN_T  _ZN4ListIP6WidgetE9add_frontES1_ strtold _GLIBCXX_HAVE_CEILL 1 _GLIBCXX_HAVE_FLOAT_H 1 _GLIBCXX_HAVE_LIMIT_VMEM 0 _GLIBCXX98_USE_C99_MATH 1 SYS_CREATE_WINDOW 22 _GLIBCXX_INCLUDE_NEXT_C_HEADERS  _GLIBCXX_HAVE_SQRTL 1 _GLIBCXX_HAVE_FCNTL_H 1 __DBL_MIN__ double(2.22507385850720138309023271733240406e-308L) __cpp_rvalue_references 200610 KEYQUEUE_SIZE 16 __GNUG__ 8 _GLIBCXX_HAVE_ETIME 1 _ZN10win_info_tC4Ev _GLIBCXX_END_NAMESPACE_CXX11 } _GLIBCXX_HAVE_FLOORL 1 _GLIBCXX_HAVE_EPERM 1 strtod __glibcxx_assert(_Condition)  SYS_SEND_MESSAGE 28 strtol SYS_UPDATE_WINDOW 26 SYS_EXIT 1 _GLIBCXX_PACKAGE_BUGREPORT "" _GLIBCXX_HAVE_ENOSPC 1 uint64_t _GLIBCXX_STD_A std _GLIBCXX_VISIBILITY(V) __attribute__ ((__visibility__ (#V))) _GLIBCXX_END_NAMESPACE_CONTAINER  atexit _ZN4ListIP6WidgetE5clearEv _Z12CreateWindowP10win_info_t GNU C++14 8.2.0 -mtune=generic -march=x86-64 -ggdb3 -g -Os __cpp_return_type_deduction 201304 _GLIBCXX_HAVE_EXPL 1 _GLIBCXX_USE_GETTIMEOFDAY 1 SYS_UNLINK 10 SYS_DESTROY_WINDOW 23 _GLIBCXX_HAVE_WCSTOF 1 WINDOW_FLAGS_NODECORATION 0x1 __GLIBCXX__ 20180726 _GLIBCXX_HAVE_EBADMSG 1 _GLIBCXX_USE_LONG_LONG 1 _GLIBCXX_BEGIN_EXTERN_C extern "C" { _GLIBCXX_END_NAMESPACE_ALGO  _GLIBCXX98_USE_C99_WCHAR 1 __GXX_WEAK__ 1 _GLIBCXX_NOEXCEPT_IF(_COND) noexcept(_COND) get_length _GLIBCXX_HAVE_UNISTD_H 1 srand __cpp_unicode_characters 200704 _GLIBCXX_HAVE_CEILF 1 _GLIBCXX_HAVE_SYS_STAT_H 1 KEY_F8 263 _GLIBCXX_BEGIN_NAMESPACE_CXX11 namespace __cxx11 { __cpp_binary_literals 201304 widgets __STDC_LIMIT_MACROS  _GLIBCXX_USE_C99_CTYPE_TR1 1 _GLIBCXX_HAVE_STRERROR_R 1 convertToDoomKey KEY_F10 265 __cpp_init_captures 201304 mbstowcs DESKTOP_SUBEVENT_WINDOW_DESTROYED 1 _GLIBCXX_HAVE_EOWNERDEAD 1 _Z16memcpy_optimizedPvS_m SYS_TIME 13 SYS_RECEIVE_MESSAGE 29 _GLIBCXX_HAVE_FABSF 1 _GLIBCXX_HAVE_SINCOSL 1 _GLIBCXX_MANGLE_SIZE_T m _GLIBCXX_HAVE_SYS_IPC_H 1 _GLIBCXX_HAVE_STDLIB_H 1 KEY_F7 262 _GLIBCXX_HAVE_INT64_T_LONG 1 __EXCEPTIONS 1 _GLIBCXX_USE_WEAK_REF __GXX_WEAK__ List<Widget*> SYS_LINK 9 _GLIBCXX_RELEASE 8 _GLIBCXX_HAVE_GETIPINFO 1 _GLIBCXX_USE_C99_STDLIB _GLIBCXX11_USE_C99_STDLIB _GLIBCXX_HAVE_LIMIT_RSS 1 _ZN4ListIP6WidgetE10get_lengthEv at_quick_exit _GLIBCXX_ATOMIC_BUILTINS 1 _GLIBCXX_HAVE_STRING_H 1 _GLIBCXX_USE_NOEXCEPT noexcept _GLIBCXX_PACKAGE__GLIBCXX_VERSION "version-unused" _GLIBCXX_HAVE_FREXPF 1 _GLIBCXX_HAVE_EIDRM 1 KEY_STATE_CAPS 1 DESKTOP_SUBEVENT_WINDOW_CREATED 2 _GLIBCXX_HAVE_ACOSF 1 _GLIBCXX_RES_LIMITS 1 _GLIBCXX_USE_C99_MATH_TR1 1 _STDDEF_H_  _GLIBCXX_HAVE_USLEEP 1 WINDOW_EVENT_KEYRELEASED 4 __cpp_runtime_arrays 198712 _GLIBCXX11_USE_C99_WCHAR 1 lldiv _GLIBCXX_HAVE_SINL 1 _GLIBCXX_HAVE_ISWBLANK 1 _ZN4ListIP6WidgetE10replace_atEjS1_ _GLIBCXX_USE_C99_FENV_TR1 1 GNU C++14 8.2.0 -m64 -mtune=generic -march=x86-64 -g -O0 -std=c++14 -fno-exceptions -fPIC _Z11SendMessagem13ipc_message_t uintptr_t /mnt/e/OneDrive/Lemon/LibLemon/build SendMessage queue_size ../src/ipc.cpp __mlibc_uintptr DrawBitmapImage _Z10surfacecpyP7SurfaceS0_8Vector2i _Z8DrawRectiiii10RGBAColourP7Surface _Z15DrawBitmapImageiiiiPhP7Surface bmp_buffer_offset fb_info_t size_aligned PointInRect rect_t bmpHeader _Z10surfacecpyP7SurfaceS0_8Vector2i4Rect colour_i memset64_optimized _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface memset32_optimized _Z11PointInRect4Rect8Vector2i srcBuffer DrawRect 20bitmap_file_header_t surfacecpyTransparent srcRegion _Z12DrawGradientiiii10RGBAColourS_P7Surface FBInfo _Z18memset32_optimizedPvjm _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i address srcHeight fbInfo DrawGradient bmpBpp rowSize _Z8DrawRect4Rect10RGBAColourP7Surface pixelSize magic CreateFramebufferSurface surfacecpy _Z24CreateFramebufferSurface6FBInfoPv bmp_offset _Z20DrawGradientVertical4Rect10RGBAColourS0_P7Surface _Z18memset64_optimizedPvmm _Z5floord _Z8DrawRectiiiihhhP7Surface destBuffer ../src/gfx/graphics.cpp srcWidth colour DrawGradientVertical yOffset overflow _ZN4ListIP6WidgetEC2Ev _ZN6WindowD2Ev _Z11PaintWindowP6Window HandleMouseUp __in_chrg _Z15HandleMouseDownP6Window8Vector2i _Z13HandleMouseUpP6Window8Vector2i ListNode _PaintWindow AddWidget ../src/gfx/window/window.cpp _ZN8ListNodeIP6WidgetEC2Ev _Z19HandleMouseMovementP6Window8Vector2i wininfo _Z12_PaintWindowPvi widget _ZN4ListIP6WidgetED2Ev _Z13_CreateWindowP10win_info_t _CreateWindow HandleMouseMovement ~Window _Z14_DestroyWindowPv widgetBounds _ZN6WindowC2Ev current _ZN6WindowD4Ev HandleMouseDown _DestroyWindow _Z9AddWidgetP6WidgetP6Window _ZN8ListNodeIP6WidgetEC4Ev _ZN6WindowC4Ev _Z13_CreateWindowP10win_info_tPPvS2_ _Znwm operator delete [] _Znam operator delete _ZdlPv _ZdaPv _ZdaPvm _ZdlPvm operator new operator new [] ../src/runtime.cpp     �@     �@      U�@     @      �U�                    �@     �@      T�@     @      �T�                 �      �       0�                                 P      Q       S                                 v p @&��e     �"�              v p ��e     �"�                 �      Q       5�                 �      Q       6�                      Z      c       Uc      �       \�      �       �U�                    Z      c       Tc      �       �T�                       Z      c       0�c      �       V�      �       v��      �       V                  }      �       S                    �      �       U�      �       �U�                    �      �       T�      �       ��                      �      �       Q�      |       V|      �       �Q�                      �      �       R�      ~       \~      �       �R�                      �      �       X�      �       _�      �       �X�                      �      �       Y�      �       ^�      �       �Y�                       �      �       0��      _       ]_      q       }�q      �       ]                            9       U9      �       V�      �       �U�                            <       T<      �       ]�      �       �T�                                  Q       �       �Q�                    a      �       \�      �       �U                       0      3       0�3             S             s�             S                    a      �       U�      -       V-      0       �U�                       �      �       S�      �       �X�      �       s���|��      �       S                                     S       $       �T$      %       s���|�%      ,       S                      q      �       R�      �       S�      �       R�             S                    �      �       R�      �       \�             R      /       \                    A      M       UM      a       �U�                            A      I       TI      Z       SZ      ^       T^      _       �T�_      `       S`      a       �T�                      )      u       Uu      �       �U��      A       U                      )      z       Tz      �       �T��      A       T                 �      A       X                 �      A       R                  �      �       Q                 �      A       [                 �      A       Z                  �      ;       S                  �      <       V                    �              P      :       Q                          S      �       U�      �       �U��      �       U�      �       \�      )       �U�                          S      �       T�      �       �T��      �       T�      !       V!      )       �T�                           S      z       0�z      �       S�      �       S�      �       0��      �       T�      �       0��      !       T                           S      �       0��      �       P�      �       P�      �       0��      �       S�      �       0��      !       S                  
             U                          *      *       R��*      1       R�0��V      V       R��V      [       R�x���      �       �P��      �       y��P��      �       �P��      �       0��P��             R�P�                                                       p r �              P       *       v�r �*      1      
 v�v ��>      J       v�r �J      P       PP      V       v�r �V      [      
 v�v ��i      |       v�r �|             Q      �       R�      �      
 v�v ���      �       v�q ��      �       ]                                      $       | v��$      1       \;      H       | v��H      [       \i      t       v�| �t      w       Pw      �       v�| ��      �       v�| �                    7      M       UM      S       P                                                              '      U       UU      j       Vj      �       U�      �       V�      �       U�      �       V�      �       U�      �       V�             U      /       V/      �       U�      �       V�      �       U�      �       V�      �       U�      �       V�      ~	       U~	      �	       V�	      �	       U�	      �	       V�	      v
       Uv
      }
       V}
      ~
       �U�                         '      e       0�e      j       1�j      r       0�r      �	       1��	      �	       S�	      x
       0�x
      |
       S|
      ~
       P                                                  u      �       P�      �       P�      �       P�      !       P/      �       P�      �       P�      �       u�      �       u�      �       P�      	       u	      +	       P+	      Y	       uY	      t	       Pt	      ~	       u~	      �	       v�	      �	       P
      v
       P                     �      �       0��      �       P�      �       p�                         �      �       0��      �       S�      �       R�      �       s��      �       S                     M      T       0�T      �       S�      �       s�                       �      �       0��      �       Q�      �       q��      �       p�                       z      }       0�}      �       P�      �       p��      �       P                          %       P%      6       S                  &      C       P                            .        U.       ^        �U�                              ,        T,       ]        \]       ^        �T�                         V        S                                   v u��       W        V                 �      �       	��                  "      B       X                 Z       `        R                     �      �       0��      �       P�      �       P                     j      q       0�q      �       P�      �       P                     E      G       0�G      Z       P[      i       P                      �      �       U�      D       ]D      E       �U�                    �      �       P�      B       \B      E       P                   �      �       0��             S      "       s�"      ?       S                               P                    %      D       UD      �       ��                      %      1       T1      �       ^�      �       �T�                            j      y       Py      �       ]�      �       \�      �       ]�      �       0��      �       ]�      �       0�                  _      �       S                    I      f       P�      �       P                    �      �       \�      �       |��      �       \                ~      �       ��                  ~      �       ]�      �       \                 �      �       0�                  �      �       9��      �       V                  �      �       P                  �      �       ^                  �      �       ��                  �      �       V                   �      �       0��      �       ]                 �      �       0�                             @       ]@      B       s �PB     "B      t       ]t      �       s �PB     "                       �       V                     t      ~       P~      �       T�      �       ]                                   U      $       S$      %       �U�                        #       P                 K       m       
 �XB     �                                  U                                  T                         .        Q                      &       ;        U;       ?        r y "�J       K        U                            n               U       �        V�       �        \�       �        �U��              \             �U�                        �       �        V�       �        \�       �        �U��              \                    �       �        P�              V                           �       �        0��       �        S�       �        V�       �        S�       �        V             S                  @      �       _                  �      �       \�      b       \                        �      �       P�      �       V�      �       P�      @       V                       �      �       p } ��      �       v } ��      �       p } ��      @       v } �                          �             S      2       p�2      �       | P-f     �\-f     ���      �       S�      �       | P-f     �\-f     ��                                       R             R      �       S�      �       | P-f     �\-f     ���      _       S                    @      �       V      ]       V                 �      �       V                   �      �       q ����4$v "��      �       q����4$v "�                   �      �       0��      �       Q                                           0�             1�             2�      &       3�&      0       4�0      :       5�:      D       6�D      N       7�                 �      �       \                     <      O       QO      R       q�]      c       Q                     ,      F       	��F      O       QO      ]       	��]      c       Q                 �      �       \                                      0�               P       %        0�0       ?        P                         (        Q                            �       U�      �       S�      �       �U�                      �      �       U�      �       �U��      0       U                      �      �       T�      �       �T��      0       T                    �             R             r�                    O       W        PW       n        R                      �       �        s v ��       �        P�       :       s v �                    T      h       Ph      �      	 X-f                             \      |       R|      ~       S~      �       R�      �       0��      �       S                    |      ~       0��      �       0��      �       V                                                        .      _       P�      �       P�      �       P�      �       s��             P2      D       P}      �       P�      �       P�      �       P�      �       P�      
       p~�      "       p~�6      p       Pq      �       P�      �       P�      �       P�      �       P�      �       P�      �       P�      �       P                     6      `       ȟ`      m       Ps      �       S                 L      c       S                        ~      �       P�      �       v��      �       PT      �       v�                       �      �       S�      �       \T      ^       S^      c       \                        1      @       ��}�@      D       TD      M       ��}�M      Q       UQ      R       ��}�                 R      R       P                 8
      C
       0�                  �      �       P                    �      V	       SV	      ]	       T                               �      �       0��      �       1��      �       2��      �       1�	      	       3�	      *	       0�*	      ;	       1�;	      L	       2�L	      ^	       3�                       �      �       S�      �       R�      �       s��      �       S                      �       �        P�       �        S�       �        P                  h       o        P                    
             P      S       V                                 Y      S       �\                  �      !       S!      S       V                  �      �       V                    ?      C       PC      S       \                     P      h       1�h      �       S�      �       S                           �       0��             T$      0       0�                    t	      x	       p  $0*��x	      6
       s  $0*��                    y	      �	       p  $0*���	      5
       p  $0*��                          )       U)      *       �U�                    �       �        U�       �        U                 �       �        0�                      �       �        U�       �        Z�       �        U                      �       �        T�       �        [�       �        T                     �       �        1��       �        Y�       �        Q                        '       8        R8       @        r�@       L        RS       �        R                    [       q        X�       �        X                                 0�                   �      =       ���=      A       U                 F             ���                        �      �       0��      �       1��             2�             3�                    �       _       ���_      h       U                                      U       �        V�       �        �U�                                      T       �        \�       �        �T�                                 0�                  c       �        S                  �
      �
       U                   N	      v	       �6f     ��	�#��v	      �	       p  $
@ $-( �                         v	      �	       0��	      �	       \�	      �	       U�	      �	       |��	      m
       \                    3	      7	       P7	      

       S                    I	      M	       PM	      k
       V                       �	      �	       p�v�15�1� ��	      
       �6f     �
��15�1� �
      
       P
      e
       S                    �      �       T�      	       �T�                  �      �       Q�      	       �Q�                  �      	       T                   �      �       t��      �       t q "#��      �       t q "#��      	       t q "#�                     �      �       P�      �      
 q 
@p "��      	      
 q
@p "�	      	      
 q 
@p "�                 �      	       r u "�                   �      �       t����      �      
 q  x �"�	      	      
 q  x �"�                  �      �       Q                  �      �       P                     �      �       p�0$0&��      �       U�      �       p�0$0&�                    �      �       s ���      �       s ��                    �      �       P�      �       P                      �      �       U�      �       V�      .       �U�                       �      �       U�      �       \�      �       V�      �       \�      +       V                           �      �       U�      �       U�      �       P�      �       U�             P
      #       P                    �      �       S�      *       S                        )       \                     �      �       0��      �       S�      �       S                        z       P                        4      E       QE      O       UO      O       q@�O      r       Qr      z       x�}�                  4      >       0�                       *       0�                      �      �       q �0$0&��      �       S�      �       q �0$0&�                      �      �       pv3��      �       p 3��      �       �6f     �:3�                   {      �      	 �6f     �             ]                      �      �       S�      �       U�      �       P                     {      �       :��      �       ^�      �       :��      �       ^�             S                   {      �       :��             \                      �      �       U�      �       �U��      �       U                       �      Y       PY      g       p��g      	       P             P                      �      s       Us             �U�      �       U                          s       Us             �U�                    �      �       U�      J       �U�                    �      �       T�      J       �T�                    �      �       Q�      J       �Q�                      �      �       R�      E       VE      J       �R�                      �      �       X�      G       \G      J       �X�                      �      �       Y�      I       ]I      J       �Y�                        5       P                      W      n       Un      �       S�      �       �U�                      W      f       Tf      �       V�      �       �T�                      W      ^       Q^      �       \�      �       �Q�                    W      z       Rz      �       �\                    2      ?       U?      W       �U�                    2      :       T:      W       �T�                    2      5       Q5      W       �Q�                    2      C       RC      W       �R�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                    �      �       Q�      �       �Q�                      a       �        U�       �        [�       �       U                    a       {        Q{       �       \                    �       �       Z�      �       z�                              $       S$      3       s p �<      A       s p �P      b       t r �b      h       t z 2$q "��                    �       �        S�       ~       S                        $       0�P      h       0�                                    $       Y$      +       p 1$y "�+      3      
 p 1$y "#�3      <      
 p1$y "#�<      A       p 1$y "�P      h       Ph      m       r 1$p "�m      u      
 r 1$p "#�u      ~      
 r1$p "#�                            >       r u z " $ &1$`�e     "�>      H      # z 2$q "�u z " $ &1$`�e     "�P      b       r u z " $ &1$`�e     "�b      ~      # z 2$q "�u z " $ &1$`�e     "�                       a       �        1��       �        P�       �        0��       �        P�      �       P                      X      i       Ui      /       V/      2       �U�                        X      u       Tu      �       S�      �       Q�      2       �T�                    X      v       Qv      2       �Q�                  )      +       s�                  �             p 31�                                    U       ^        �U�                                    T       ^        �T�                                         0�       4        P:       B        PU       ]        P]       ^        p 1'�                      
               Y       U        y x "�U       X        y x "#�X       ^        y x "�                                     Z       U        z x "�U       X        z x "#�X       ^        z x "�                    0       :        R>       U        R                    �      �       U�      �       �U�                    �      �       T�      �       �T�                      �      �       U�      O       VO      X       �U�                        �      �       T�      �       R�      Q       \Q      X       �T�                      �      �       Q�      S       ]S      X       �Q�                           -       U6      >       U                       �      	       0�	      6       T6      9       t�>      G       T                    �      M       PM      W       U                  �s@     �s@      P                       �s@     �s@      t �4�-�-  Bp �4�-��s@     �s@      t �4�-�-  Bq �4�-��s@     �s@      a�s@     �s@      t �4�-�-  Bq �4�-�                    �s@     �s@      P�s@     �s@      Q                      Is@     Rs@      URs@     _s@      S_s@     �s@     	 �;f                       r@     +s@      S                     �r@     �r@      0��r@     �r@      P�r@     �r@      p�                  .r@     ,s@      V                  >r@     >s@      \                  �q@     r@      S                 �q@     r@     
 ��B     �                �q@     �q@      S                   q@     q@      0�q@     'q@      P                  �n@     o@      U                    "o@     Jo@      SJo@     No@      T                  ^o@     to@      P                   Oo@     {o@      @=$�{o@     �o@      S                            fu@     �u@      U�u@     .v@      \.v@     7v@      �U�7v@     �v@      \�v@     �v@      U�v@     �v@      �U�                    �u@     6v@      P7v@     Vv@      P                  Av@     �v@      S                      nv@     �v@      P�v@     �v@      V�v@     �v@     	 P9f                       tv@     �v@      ]                      Lv@     Rv@      ^Rv@     Vv@      UVv@     �v@      ^                      �t@     �t@      U�t@     �t@      �U��t@     fu@      U                        �k@     �k@      U�k@     �k@      \�k@     �m@      ]�m@     �m@      �U4�U $@N$,( �                              �k@     �k@      T�k@     l@      Sl@     l@      �T�l@     $l@      S$l@     5l@      �T�5l@     �m@      S�m@     �m@     	 9f                             �k@     �k@      Q�k@     Rl@      VRl@     Tl@      �Q�Tl@     �m@      V                  �m@     �m@      U                           m@     m@      0�m@     !m@      1�!m@     +m@      2�+m@     5m@      3�5m@     �m@      4�                    �j@     �j@      P�j@     �k@      \                    �j@     �j@      P�j@     �k@      V                     qj@     �j@      0��j@     �j@      P�j@     �k@      S                      Oj@     `j@      U`j@     dj@     	  �e     dj@     qj@      �U�                    Oj@     dj@      Tdj@     qj@      �T�                      0j@     >j@      U>j@     Bj@      TBj@     Oj@      �U�                              -g@     @g@      X@g@     Cg@      x��g@     �g@      0��g@     �g@      1��g@     �g@      2��g@     �g@      3�*i@     /i@      0�/i@     =i@      R                          ee@     �e@      U�e@     �e@      S�e@     �e@      s��e@     �e@      S�e@     �e@      �U�                  �e@     �e@      Q                      �e@     �e@      D} ��e@     �e@      E} ��e@     �e@      D} �                    �e@     �e@      T�e@     �e@      \                          �c@     �c@      U�c@     �c@      ]�c@     �c@      U�c@     5d@      ]5d@     ee@      �U�                          �c@     �c@      T�c@     �c@      �T��c@     �c@      T�c@     Xe@      \Xe@     ee@      �T�                  �c@     Xe@      S                  �c@     Xe@      V                    ed@     kd@      Pkd@     Xe@      ]                  4e@     We@      P                    �c@     �c@      P�c@     �c@      p�                             �d@     �d@      U�d@     �d@      U�d@     �d@      U�d@     �d@      Ue@     
e@      Ue@     e@      0�e@     )e@      U                             �d@     �d@      T�d@     �d@      T�d@     �d@      T�d@     �d@      Te@     
e@      Te@     e@      0�e@     !e@      T                                      zd@     �d@      T�d@     �d@      p 0$0&:$��d@     �d@      T�d@     �d@      p 0$0&:$��d@     �d@      T�d@     �d@      p 0$0&:$��d@     �d@      T�d@     �d@      p 0$0&:$��d@     e@      Te@     
e@      |�r 0$0&:$�
e@     e@      T                    �b@     �b@      U�b@     �c@      �U�                 �b@     �c@      Q                   �c@     �c@      0��c@     �c@      1��c@     �c@      2��c@     �c@      3��c@     �c@      4�                  �b@     �c@      a�                   �b@     �b@      u  $ &
H�<f     "�b@     �b@      �U $ &
H�<f     "                    �b@     �b@      u  $ &
H�<f     "�b@     �b@      �U $ &
H�<f     "                  �b@     �c@      Z                    ob@     �b@      U�b@     �b@      �U�                   ob@     �b@      u  $ &
H�;f     "��b@     �b@      �U $ &
H�;f     "�                    �c@     �c@      U�c@     �c@      �U�                            �v@     �v@      0��v@     �v@      S�v@     �v@      s�zw@     }w@      0�}w@     �x@      S�x@     �x@      s��x@     [y@      S[y@     ^y@      s�                            zw@     }w@      Q}w@     �y@      \�y@     �y@      \�y@     �y@      \�y@     �y@      \�y@     �y@      \                  �w@     �x@      ]                      �_@     �_@      U�_@     mb@      Smb@     ob@      �U�                  <a@     �a@      [                     <a@     Ya@      0�Ya@     �a@      R�a@     �a@      r�                  ta@     �a@      Z                  �a@     Kb@      Z                     �a@     �a@      0��a@     7b@      R7b@     :b@      r�                    b@     Nb@      p ��Nb@     fb@      r2$D�e     "���                 k^@     r^@      0�                  7^@     ;^@      U                      �W@     _X@      U_X@     �]@      S�]@     �]@      �U�                    �W@     mX@      TmX@     �]@      �T�                         �[@     �[@      r  $ &3$$�B     "�[@     �[@      P�[@     �[@      Q�[@     �[@      p��[@     �[@      q�                  X@     �]@      ^                  �\@     ]@      Q                  KX@     �]@      ]                      �X@     �X@      P�X@     Y@      PY@     (Y@      P                     KX@     KY@      0�KY@     p]@      \p]@     �]@      Q                         KX@     �X@      0��X@     �X@      V�X@     ,Y@      0�,Y@     {]@      V{]@     �]@      P                     �[@     �[@      p 3$��B     "�[@     �[@      p 3$��B     "�[@     �[@      p3$��B     "                    �]@     �]@      P�]@     �]@      ��e     �s�"�                �Z@     �[@      Y                  �Z@     )[@      Q                                  �Z@     �Z@      0��Z@     �Z@      P�Z@     �Z@      p��Z@     �Z@      x�)[@     )[@      R)[@     -[@      y r "�-[@     5[@      P5[@     8[@      pw�8[@     ;[@      y r "�;[@     S[@      QS[@     �[@      R                  G[@     �[@      P                   �W@     �W@      0��W@     �W@      1��W@     �W@      2��W@     �W@      3�                     �W@     �W@      0��W@     �W@      u �W@     �W@      P�W@     �W@      u�p "��W@     �W@      P                                �e@     Cf@      UCf@     Df@      �U�Df@     [f@      U[f@     ~f@      S~f@     �f@      s��f@     �f@      �U��f@     �f@      S�f@     �f@      �U�                          Jf@     ~f@      S~f@     �f@      s��f@     �f@      �U��f@     �f@      S�f@     �f@      �U�                      `f@     �f@      \�f@     �f@      |��f@     �f@      |�                  !n@     nn@      S                      v      �       U�      �       S�      �       �U�                      b      t       Ut      u       �U�u      v       U                     b      t       Ut      u       �U�u      v       U                      #      +       U+      a       Sa      b       �U�                            #      /       T/      0       �T�0      B       PB      E       TE      P       PX      ]       P                                  U      #       R                                T      #       X                 �      �       U                    �      �       U�      �       R                 �      �       X                 �      �       R                 �      �       Q                 �      �       T                 �      �       U                 �      �       U                      :      B       UB      �       S�      �       �U�                     :      B       0�B      r       V|      �       V                      �             U      9       V9      :       �U�                            (       S(      4       s�4      8       S                               	 v��s �      ,       U                   !      ,       u  $ &pv "�/      3       U                    �      �       U�      �       X                    �      �       T�      �       Z                    �      �       Q�      �       Y                     �      �       0��      �       P�      �       P                   h      v       u�� $ &pu "�v      �       P                  �             U      F       �U�                         .       Z.      C       z�C      F       Z                 ?      C       u�                 ?      C       u�                 ?      C       [                 ?      C       u�                      /      B       UB      �       S�      �       �U�                  |      �       ]                 |      �       V                 |      �       \                                 �        U�              S      &       �U�&      '       S'      /       �U�                                 �        T�              \      &       �T�&      *       \*      /       �T�                         �       �        0��       �        ]�       �        }��              ]&      ,       ]                      �       �        q �0$0&��       �        ^�       �        q �0$0&�                         �       �        V�       �        U�              V      %       U&      (       V                    �       �        P�       �        P                 )       1        U                                b      �       U�             �U�      (       U(      �       �U��             U      k       �U�k      s       Us      �       �U�                            '       T'      )       t�)      O       T                                 b      �       0��      �       1��      �       0��             1�      h       0�h      ~       1�~      f       0�f      k       1�k      ~       0�~      �       P�      �       S                                 P      S       Rn      �       V                         b      b       0�b      b       1�b      b       2�b      b       3�b      �       4�      9       4�9      �       S�      �       s��      �       4�                
b      b       0�                  [      a       P                          �       S�      �       s�                  a      ~       P                  ,      �       \                    J      L       Si      �       S                                     0�       7        S7       :        s�                                   !�               s!�       :        s"�                       �       �        S�       �        R�       �        s��       �        S                    �             U             u{�      %       U                    �      
       T
             t�      %       T                      �      �       U�      �       p 2$u "��      �      
 p 2$u "#��      �      
 p2$u "#�                      �      �       T�      �       t p "��      �       p t "#��      �       p t "�                      �      �       Q�      �       q p "��      �       p q "#��      �       p q "�                   �      �       0��      �       P�      �       p�                  �      �       x ��                      �      �       U�      �       p 2$u "��      �      
 p 2$u "#��      �      
 p2$u "#�                      �      �       T�      �       t p "��      �       p t "#��      �       p t "�                   �      �       0��      �       P�      �       p�                    l      �       U�      �       u}��      �       U                     l      o       To      |       t x "�|      �       t x "1�                     l      o       Qo      |       q x "�|      �       q x "1�                   l      o       0�o      |       X                  �      �       p ��                    K      T       UT      c       u}�c      l       U                     K      M       TM      `       t p "�`      c       p t "1�                   K      M       0�M      `       P                                   U      ?       p 1$u "�?      B      
 p 1$u "#�B      K      
 p1$u "#�                                   T      ?       t p "�?      B       p t "#�B      K       p t "�                                   Q      ?       q p "�?      B       p q "#�B      K       p q "�                                0�      ?       P?      B       p�                  6      K       x ��                                   U             p 1$u "�            
 p 1$u "#�            
 p1$u "#�                                   T             t p "�             p t "#�             p t "�                                0�             P             p�                      �      �       U�      �       u x "��      �       u x "#��             u x "�                      �      �       T�      �       t x "��      �       t x "#��             t x "�                      �      �       Q�      �       q x "��      �       q x "#��             q x "�                   �      �       0��      �       X�      �       x�                      f      q       Uq      �       S�      �       �U�                      �      �       U�      �       S�      �      	 ��
 �                      �      �       T�      �       V�      �       �T�                        �      �       P�      �       \�      �       ]�      �       P                 �      �       0�                      �      �       0��      �       { | ��      �       { | #�                    �      �       P�      �       ��                                 P      �       ��                 

 3      3       P3      �       ��                   �      �       U�      �       u}�                   �      �       T�      �       t}�                

 3      3       P3      �       ��                 3      �       ��                 3      �       ��                 3      �       S                   3      �       X�      �       x}�                

 3      3       0�3      �       ^                	

   3      3       ����3             _�      �       _                    r      u       p y "�u      �       P                
 3      �       Q                    F      �       U�      �       �U�                  F      �       T�      �       �T�                    F      u       Ru      �       �D                  �      �       Y                   �      �       X�      �       Z�      �       Z                    �      �       ]�      �       [�      �       [                        �      �       ^�      �       S�      �       S�      �       ~ u "��      �               � $ &1$x "u "�                      �      �       S�      �       V�      �       V�      �       ��u "�                      �      �       R�      �       \�      �       \�      �       ��u "�                   �      �      
 �Ur "y ��      �      
 �Ur "y �                 �      �       T                    L      �       p 5��      �               �5�                    �      �       z p "��             z p "#�             z p "#�             z p "#�             z p "#�      �       z p "#��      �       z p "�                    �             { p "�      "       { p "#�"      +       { p "#�+      0       { p "#�0      9       { p "#�9      �       { p "#��      �       { p "�                    �      >       s p "�>      F       s p "#�F      K       s p "#�K      T       s p "#�T      Y       s p "#�Y      �       s p "#��      �       s p "�                    �      b       v p "�b      g       v p "#�g      p       v p "#�p      u       v p "#�u      ~       v p "#�~      �       v p "#��      �       v p "�                    �      �       | p "��      �       | p "#��      �       | p "#��      �       | p "#��      �       | p "#��      �       | p "#��      �       | p "�                    �      �       R�      �       r��      �       R                  N      �       T�      F       �T�                  ~      F       X                  �      F       Y                  �      F       [                  �      =       S                  �      F       Z                        �      �       u p "��      �       \�             u p "�              p u "#�"      <       \                 �      F       T                    j      �       P�      C       VC      F               �2$�                      �      �       p 2$y "��      �      
 p 2$y "#��      �      
 p 2$y "#��      �      
 p 2$y "#��             
 p 2$y "#�       "      
 p2$y "#�"      %       p 2$y "�                      �      �       p 2${ "��      �      
 p 2${ "#��      �      
 p 2${ "#��      �      
 p 2${ "#��             
 p 2${ "#�       "      
 p2${ "#�"      (       p 2${ "�                      �      �       p 2$s "��      �      
 p 2$s "#��      �      
 p 2$s "#��      �      
 p 2$s "#��             
 p 2$s "#�       "      
 p2$s "#�"      +       p 2$s "�                      �             p 2$z "�      
      
 p 2$z "#�
            
 p 2$z "#�            
 p 2$z "#�             
 p 2$z "#�       "      
 p2$z "#�"      .       p 2$z "�                      �             x p "�              x p "#�       5       x p "�5      <      
 x p "
@�                    �       �        U�       N       �U�                  �       �        T�       N       �T�                  �       N       [                  �       J       P                  �       E       S                  �       N       X                   �       �       
 �Uz "{ �$      :      
 �Uz "{ �                 �       N       T                    �       �        Y�       K       VK      N               �3�                    �       �        p y "��       �        p y "#��       �        p y "#��       (       p y "#�(      -       p y "�                    �       �        s y "��               s y "#�       	       s y "#�	      (       s y "#�(      0       s y "�                    �              x y "�             x y "#�             x y "#�      (       x y "#�(      3       x y "�                    �       �        Z�       $       z�$      D       Z                            F        TF       �        �T�                  (       �        X                      8       D        PD       E       %         �t u "1$ $ &        "�E       �        P                  ;       �        Y                          I       M        u z "�M       U        SU       k        u z "�k       n        u z "#�p       �        S�       �        u z "�                     ;       r        Tr               t�       �        T                           F        ZF       �        [                      I       Q        z 1$p "�Q       Y       
 z 1$p "#�Y       n       
 z 1$p "#�n       p       
 z1$p "#�p       u        z 1$p "�                      I       ^        z 1$y "�^       f       
 z 1$y "#�f       n       
 z 1$y "#�n       p       
 z1$y "#�p       x        z 1$y "�                      I       k        x z "�k       n        x z "#�n               x z "�       �       
 x z "
@�                  %      `       U`      �       �U�                  %      `       T`      �       �T�                    %      .       Q.      �       �Q�                  %      `       R`      �       Z                  S      �       P                     `      q       Xq      s       Us      �       X                 `      �       Y                  .      �       Q                  �      �       U                      �             T             �T�             T                      �             Q             �Q�             Q                      �      �       R�             �R�             R                  �             0�                  �             
@�                  �             ȟ                                
      [       S[      b       Qb      m       Tm      z       ]z      �       Q�      �       T�      �       s�x��      �       Q�      �       T�      �       Q�      �       T�      �       S�             t��                     
      5       R5      �       Z�             R                 
             0�                               U                            Q       TQ      �	       �T��	      �	       T                            Q       QQ      �	       �Q��	      �	       Q                            ;       R;      �	       �R��	      �	       R                  2      �	       0�                  2      �	       
@�                  2      �	       ȟ                              J      �       S�      �       T�      �       s���      �       Q�      	       T	      	       Q	      I	       TI	      M	       ]M	      T	       QT	      u	       Tu	      	       S	      �	       t��                     J      u       Ru      M	       ZM	      �	       R                 J      Q       0�                  �	      �	       U                      �	      �	       T�	      R       �T�R      V       T                      �	      �	       Q�	      R       �Q�R      V       Q                      �	      �	       R�	      R       �R�R      V       R                  �	      R       0�                  �	      R       
@�                  �	      R       ȟ                                �	      3
       S3
      f
       Tf
      s
       ]s
      �
       Q�
      �
       T�
      �
       s���
      �
       Q�
      	       T	             ]             Q      9       T9      C       SC      R       t��                     �	      �	       R�	             Z      R       R                 �	      �	       0�                  V      Z       U                      V      �       T�      "       �T�"      &       T                      V      �       Q�      "       �Q�"      &       Q                      V      �       R�      "       �R�"      &       R                  x      "       0�                  x      "       
@�                  x      "       ȟ                          �       P�             y�}�              P                  �      "       T                 �      �       0�                    �      �       P�             p{�             P                      �      �       T�      �       R�      �       r��      �       r}��             R                    �      �       0��      �      	 p y #��                  &      *       U                      &      ~       T~      ^       �T�^      b       T                      &      ~       Q~      ^       �Q�^      b       Q                      &      ~       R~      ^       �R�^      b       R                  H      ^       0�                  H      ^       
@�                  H      ^       ȟ                    O      �       P�      K       v�}�K      Z       P                  V      ^       X                 V      ~       0�                   ~      �       P�      ?       p{�?      H       P                      ~      �       X�      �       Q�      �       qx�7      H       Q                    �      �       R�      �       r��      �       ry�7      H       R                   �      �       0��      �      	 p v #��                                  �      �       t ���      �       qx����      �       t ���      �       qz����      �       t ���             q{���             t ��      +       q}���+      ^       t ��                  b      f       U                      b      �       T�      ^       �T�^      b       T                      b      �       Q�      ^       �Q�^      b       Q                      b      �       R�      ^       �R�^      b       R                  �      ^       0�                  �      ^       
@�                  �      ^       ȟ                    �      F       XF      I       x�}�I      ^       X                  �      ^       Q                 �      �       0�                     �      �       X�      �       U�      3       u~�3      ?       U                               �      �       Q�      �       q p "��      �       q p "#��             q p "#�             q p "#�      .       q p "#�.      7       q p "#�7      ?       q p "�                                �      �       Y�      �       y p "��      �       y p "#��             y p "#�             y p "#�      )       y p "#�)      7       y p "#�7      ?       y p "�                      �      �       Z�      �       z p "��      �       z p "#��             z p "#�             z p "#�      $       z p "#�$      7       z p "#�7      ?       z p "�                   �      �       0��      �       u x �                      �      �       t ���             q p "#���      ^       t ��                  b      f       U                      b      �       T�      �       �T��      �       T                      b      �       Q�      �       �Q��      �       Q                      b      �       R�      �       �R��      �       R                  �      �       0�                  �      �       
@�                  �      �       ȟ                    �      �       P�      �       ~�}��      �       P                  �      �       Z                 �      �       0�                   �             P      w       p{�w      �       P                      �      �       Z�             Q             qp�g      �       Q                   �      �       0��            	 p ~ #��                                  �      :       y ��:      N       qr���N      �       y ���      �       qu����      �       y ���      �       qx����             y ��      3       q{���3      �       y ��                     �      �       R�             rp�g      �       R                     �      �       T�      	       tp�g      �       T                    �      �       U�      �       u��             uq�g      �       U                  �      �       U                      �             T      �       �T��      �       T                      �             Q      �       �Q��      �       Q                      �      �       R�      �       �R��      �       R                  �      �       0�                  �      �       
@�                  �      �       ȟ                    �      �       U�      �       u�}��      �       U                  �      �       R                 �             0�                                U             u p "�      �       u p "#��      �       u p "�                                        R      2       p 2$r "�2      I      
 p 2$r "#�I      a      
 p 2$r "#�a      y      
 p 2$r "#�y      �      
 p 2$r "#��      �      
 p2$r "#�                         }       P}      �       p�                  "      �       q ��                                         X      .       p 2$x "�.      D      
 p 2$x "#�D      \      
 p 2$x "#�\      t      
 p 2$x "#�t      �      
 p 2$x "#��      �      
 p2$x "#�                                         Y      *       p 2$y "�*      ?      
 p 2$y "#�?      W      
 p 2$y "#�W      o      
 p 2$y "#�o      �      
 p 2$y "#��      �      
 p2$y "#�                                         Z      &       p 2$z "�&      :      
 p 2$z "#�:      R      
 p 2$z "#�R      j      
 p 2$z "#�j      �      
 p 2$z "#��      �      
 p2$z "#�                                 [      "       p 2${ "�"      5      
 p 2${ "#�5      M      
 p 2${ "#�M      e      
 p 2${ "#�e      �      
 p 2${ "#��      �      
 p2${ "#�                  �      �       U                      �      �       T�      �       �T��      �       T                      �      �       Q�      �       �Q��      �       Q                      �      �       R�      �       �R��      �       R                  �      �       0�                  �      �       
@�                  �      �       ȟ                            �      <       V<      _       T_      b       v�v�b      s       Qs      v       v�x�v      �       Q�      �       T�      �       \�      �       V�      �       |���      �       q��                           �             P      �       Z�      �       P�      �       U�      �       z { "��      �       P�      �      	 z { "{ "�                 �      �       0�                        �      �       U�             S             �U�             U                      �      �       U�             S             �U�                              3       U3      W       SW      c       �U�c      d       U                      .      3       U3      W       SW      c       �U�                  d      h       U                      d      �       T�      M       �T�M      Q       T                      d      �       Q�      M       �Q�M      Q       Q                    d      �       R�      M       �R�M      Q       R                  �      M       0�                  �      M       
@�                  �      M       ȟ                    �      �       X�      �       x�}��             X                       �             R7      D       QD      F       UF      M       Q                      �      �       0�7      9       0�9      F      	 x 	�#�	�F      I      	 x 	�#�	�I      M      	 x	�#�	�                                   U             �U�             U                                   T             �T�             T                      �             U             �U�             U                      �      �       U�      �       �U��      �       U                      �      �       T�      �       �T��      �       T                      �      �       U�      �       �U��      �       U                      �      �       U�      �       �U��      �       U                      �      �       T�      �       �T��      �       T                      �      �       U�      �       �U��      �       U                      x      �       U�      �       �U��      �       U                      :      t       Ut      u       �U�u      x       U                      :      t       Tt      u       �T�u      x       T                        :      c       Qc      r       q  $0 $+( �r      u      & �Q�Q $�O$,(  $0 $+( �u      x       Q                        :      V       RV      l       r  $0 $+( �l      u      ' �R��R $� $,(  $0 $+( �u      x       R                            8       U8      9       �U�9      :       U                              *       T*      6       t  $0 $+( �6      9      & �T�T $�O$,(  $0 $+( �9      :       T                                     Q      1       q  $0 $+( �1      9      ' �Q��Q $� $,(  $0 $+( �9      :       Q                      �       �        U�       �        �U��       �        U                                    U       y        �U�                                   p  $0+��       x        |  $0+��                    "       &        p  $0+��&       u        s  $0+��                      '       A        p  $0+��A       p        v  $0+��p       t        p  $0+��                 T       c        �U�                 _       c        0�                 n       p        0�                      �      �       U�             S             �U�                      �      �       T�             V             �T�                      �      �       Q�      �       ^�             ^                    �      �       P�      �       \                   �      E       0�E      n       _                          �       k       Uk      r       Vr      |       U|      .       V.             �U�                  .      �       V                  L      ]       p  $0)��                T      �       \�             ��z�                �             V                     �      �       P�      �       U�             \                f      �       \�      �       ��z�                 �      �       P�      �       V                      �      �       P�      �       ]�      �       }��      �       ]�      �       }��      �       ]�      �       }�                    �      �       \�      �       |��      �       \                  �       �        S                    �       �        U�       �        �h                       t       z        0�z       �        Ks ��       �        Ls ��       �        Ks �                  /       F        U                     T       a        \a       f        |�f       o        \                  T       m        V                            "       U"      �       V�      �       �U�                       m      z       Pz      ~       T~      �       \�      �       P                 F      F       P                  -      C       P                F      m       V                    F      Y       0�Y      ^       P^      m       0�m      m       P                              	        U	       -        V-       .        p                                       T       ,        S,       .        p                         .        P                    Q       U        UU       V        �U�                  :       O        P                                   P       $        p ��e     ��$       .        P                    �      �       U�      �       �U�                        �      �       T�      �       �T��      �       T�      �       �T�                    �      �       Q�      �       �Q�                    �      �       T�      �       T                        k      x       Ux      �       S�      �       U�      �       �U�                    �       �        U�       Q       \Q      ]       �U�                    �       �        T�       ]       �T�                    �       �        Q�       Q       ]Q      ]       �Q�                    �       �        R�       Q       SQ      ]       �R�                    �       �        T�       D       VD      Q       �T} �                           )       P)      3       ^                      �       �        P�       �        S�       �        P                        -       9        U9       D        �U�D       w        Uw       �        Z                          -       =        T=       D        �T�D       Q        TQ       �        X�       �        �T�                          -       =        Q=       D        �Q�D       N        QN       i        Pi       �        �Q�                        -       =        R=       D        �R�D       W        RW       �        Y                     T       i        Pi       n        �Q�n       �        P                                      U       ,        V,       -        p                                       T       +        S+       -        p                         -        P                  x       �        P                    K       N        UN       O        �U�                    O       T        UT       _        �U�                                      U       J        ^J       K        �U�                                    T       K        �T�                                       1�"       1        S1       <        \<       ?        S                      �       �        U�       �        tD��       �        �U�                    �       �        T�       �        P                                    U       �        Q                    �      �       U�      8       �U�                            #       P#      7       S7      8       P                    �      �       U�      �       �U�                 �      �       P                    �      �       U�      �       �U�                  �      �       P                    a      f       Uf      �       �U�                  g      ~       P                    >      C       UC      a       �U�                  D      [       P                    �      �       U�      >       �U�                      �      �       T�      =       V=      >       �T�                        �      �       P�      �       S�      �       S�      5       S                 �      :       V                     �      �       S�      �       S�      5       S                                   P             s      !       Q                    �      �       U�      �       �U�                      �      �       T�      �       S�      �       p                  �      �       P                        F       R        UR       X        TX       �        V�       �        �U�                          \       m        Pm       q        Sq       �        P�       �        S�       �        P                        �       �        P             PM      f       Ps      �       P                 �       �       	 0Ge                      �       �       	 08e                                           U       A        \A       F        �U�                                      T       E        ^E       F        �T�                                     0�       "        V8       :        V                        �       �        U�       �        u~��       �        U�       �        �U�                    �       �        U�       �        u~�                      �             U      H       VH      I       �U�                         ;       SB      G       S                           B        TB       L        �T�                   <       K        u  $ &@$t  $ &�K       L        P                            
        U
               �U�                         l�@     ��@      \��@     �@      ]P�@     ��@      S��@     ��@      s���@     �@      S                 P�@     �@      V                    f�@     p�@      u�p�@     y�@      U                       �@     @�@      0���@     ��@      ~���@     ��@      VĦ@     Ȧ@      p v "1�Ȧ@     �@      V                   ��@     ��@      1���@     Ȧ@      0�                                          �@     �@      U�@     	�@      V	�@      �@      U �@     &�@      V&�@     P�@      UP�@     ~�@      V~�@     ��@      U��@     k�@      Vk�@     ��@      �U���@     ѱ@      Vѱ@     ر@      �U�ر@     ��@      V��@      �@      �U�                                                                       Z�@     f�@      U~�@     ��@      0���@     �@      U�@     +�@      UF�@     T�@      UX�@     [�@      P[�@     ��@      \��@     	�@      U�@     1�@      U7�@     `�@      Ub�@     ��@      U��@     ŭ@      Uۭ@     �@      U �@     0�@      U:�@     I�@      UX�@     b�@      Ux�@     ��@      U��@     ��@      U��@     ˮ@      U�@     *�@      U{�@     ��@      Uү@     �@      U-�@     c�@      U��@     ��@      U�@     �@      U �@     X�@      U_�@     ʱ@      Uر@     ��@      U                                     Z�@     f�@      S~�@     ��@      	����@     N�@      SN�@     ��@      	����@     ��@      S��@     ��@      	����@     |�@      S|�@     ��@      	����@     {�@      S��@     y�@      Sy�@     ��@      s��                      ��@     ��@      P��@     ʱ@      Pر@     ��@      P                  c�@     s�@      S                      H�@     [�@      U[�@     ��@      ]��@     ��@      �U�                    H�@     [�@      T[�@     ��@      �T�                    H�@     [�@      Q[�@     ��@      �Q�                      ��@     ��@      q �0$0&���@     ��@      S��@     ��@      q �0$0&�                    W�@     [�@      Q[�@     ��@      \                      d�@     s�@      Ux�@     |�@      U��@     ��@      P                       W�@     [�@      U[�@     m�@      ^m�@     s�@      ]x�@     ��@      ^��@     ��@      S��@     ��@      ^                    Z�@     [�@      T[�@     ��@      V                  �@     $�@      U                    �@     4�@      0�4�@     H�@      Q                    �@     4�@      T4�@     H�@      P                   �@     H�@      T                  ��@     Σ@      U                       ��@     ٣@      0�٣@     �@      s �U��@     �@     	 s �U#��@     
�@      s �U�                     ��@     ٣@      0�٣@     �@      V�@     �@      P                  �@     ��@      P                      �@     �@      U�@     <�@      V<�@     A�@      �U�                      �@     �@      T�@     "�@      S"�@     A�@      �T�                      ١@     �@      U�@     �@      V�@     �@      �U�                      ١@     �@      T�@     �@      S�@     �@      �T�                          �@     	�@      U	�@     �@      S�@     "�@      U"�@     ��@      sx���@     ��@      �U�                        �@     ��@      T��@     ��@      \��@     ��@      T��@     ��@      �T�                      �@     �@      Q�@     b�@      Vb�@     ��@      �Q�                      �@     �@      R�@     ��@      ^��@     ��@      �R�                            �@     	�@      U	�@     �@      S�@     "�@      U"�@     #�@      sx�#�@     #�@      S#�@     D�@      _D�@     K�@      UK�@     L�@      x�L�@     ��@      _                   #�@     5�@      ]5�@     L�@      }�L�@     ��@      ]                    ,�@     8�@      U<�@     R�@      U                  ל@     ל@      Uל@     ,�@      0�                    �@     3�@      U3�@     m�@      �U�                 7�@     7�@      R                    ��@     ϲ@      Uϲ@     ۲@      �U�                 Ѳ@     ֲ@      0�                  ��@     ��@      U��@     ��@      0�                  �@     �@      U�@     Q�@      0�                    ��@     ��@      U��@     ��@      �U�                    ��@     ��@      U��@     ��@      U                    i�@     u�@      Uy�@     ��@      U                     �@     �@      U�@     
�@      �U�                   ��@     A�@     
 �SB     �A�@     J�@      U                   ��@     A�@      
J�A�@     h�@      V                   ��@     A�@      ��A�@     g�@      S                      8�@     I�@      UI�@     j�@     	 �Df     j�@     ��@      �U�                      ��@     ��@      U��@     ş@      Sş@     Ɵ@      �U�                    �@     �@      U�@     8�@      �U�                          "�@     4�@      U4�@     f�@      Sf�@     m�@      Um�@     n�@      sx�n�@     ��@      S��@     ��@      U                          "�@     ,�@      T,�@     7�@      V7�@     ��@      vy���@     ��@      ty���@     ��@      �T�                        ��@     Ş@      PŞ@     ؞@      \؞@     �@      P�@     !�@      \                     v�@     ��@      0���@     �@      S�@     �@      s�                    ~�@     ��@      U��@     ��@      U                  ��@     ��@      0�                        ��@     �@      U�@     ��@      �U���@     ��@      U��@     ��@      �U�                      ��@     �@      U�@     ��@      �U���@     ��@      �U�                      ��@     �@      U�@     �@      �U��@     �@      U                    �@     �@      U�@     �@      �U�                      �@     7�@      U7�@     K�@      �U�K�@     L�@      U                    &�@     7�@      U7�@     K�@      �U�                      L�@     t�@      Ut�@     u�@      �U�u�@     v�@      U                    T�@     t�@      Ut�@     u�@      �U�                      Ɵ@     ՟@      U՟@     �@      �U��@     �@      U                    Ο@     ՟@      U՟@     �@      �U�                  ע@     ע@      Uע@     �@      0�                    �@     �@      U�@     �@      �U�                        m�@     ��@      U��@     ��@      �U���@     ��@      U��@     ��@      �U�                  r�@     ��@      4�                  ��@     ƥ@      P                        �@     �@      U�@     #�@      �U�#�@     )�@      U)�@     4�@      �U�                    �@     �@      U�@     #�@      �U�                          4�@     F�@      UF�@     K�@      �U�K�@     Z�@      UZ�@     e�@      �U�e�@     f�@      U                    =�@     F�@      UF�@     K�@      �U�                        
�@     %�@      U%�@     *�@      �U�*�@     ?�@      U?�@     K�@      �U�                    �@     %�@      U%�@     *�@      �U�                        K�@     _�@      U_�@     o�@      �U�o�@     ��@      U��@     ��@      �U���@     ��@      0�                    Z�@     _�@      U_�@     o�@      �U�                  ��@     ��@      U��@     ��@      0�                    X      �       U�      �       �U�                    X      �       T�      �       �T�                    X      �       Q�      �       �Q�                  �      �       P                  �             U                          �      �       P�      �       V�      �       P�             V             P                  B             S                  �      �       U                  �      �       T                  l      z       U                  l      �       T                  H      S       U                    H      k       Tk      l       �T�                    H      d       Qd      l       �Q�                    Z      g       Ug      k      ' r�Qr#����������Q#���������,( �                    G      e       Ue      �       V                  G      s       T                   G      q       Qq      �       w                       �      �       P�      C       ]C      H       P                 �      6       _                         �      �       Q�      �       P�      �       Q�      �       P�      �       V      6       V                  }      A       \                  �      �       S                   �      *       S*      -       s�-      6       S                    �      �       U�      �       S                      �      �       P�             V      	       P                  \      x       U                  \      �       T                  �      �       V                    �      �       Q�      �       S                  �      �       V                   �      �       0��      �       _                  A      E       UE      \       �U�                     E      U       SU      X       s�X      [       S                  �      �       U                            �      �       T�      7       \7      ;       Q;      <       �T�<      @       \@      A       �T�                          �             S             s v "�             s v "#�      2       s v "�2      5       t v "�<      =       s v "�                       �      �       S      2       S2      ;       T<      =       S                         �      �       0�      
       V
             v�      5       V<      >       V                      _      v       Uv      �       S�      �       �U�                        _      n       Tn      v       Qv      �       V�      �       �T�                            "       U"      (       Q(      )       �U�                      �       �        U�       X       \X      _       �U�                      �       �        T�       \       ^\      _       �T�                    �       �        P�       V       V                  5      ^       _                               P                        *      .       P.      Z       ]Z      \       ~ \      _       �T                    �       �        U�       �        �U�                      �       �        T�       �        \�       �        �T�                      �       �        Q�       �        V�       �        �Q�                    �       �        P�       �        S                  �       �        \                      H       S        US       �        S�       �        �U�                    a       e        Pe       �        \                      y       }        P}       �        V�       �        P                    
               U       H        �U�                           !        P)       9        P                            	        U	       
        �U�                      	      "       U"      1       �U�D      G       U                        	      "       T"      =       S=      D       �T�D      G       T                        	             Q      "       P"      D       �Q�D      G       Q                            "       T"      =       S=      C       �T�                          "       U"      C       �U�                    7      @       p�@      C       r  1�                        )      >       U>      V       VV      W       �U�W      X       U                        )      >       T>      U       SU      W       �T�W      X       T                      )      >       Q>      W       �Q�W      X       Q                      )      >       R>      W       �R�W      X       R                    4      >       R>      W       �R�                    4      >       Q>      W       �Q�                      4      >       T>      U       SU      W       �T�                      4      >       U>      V       VV      W       �U�                  ?      W       P                                 0�      8       R8      ;       r�                                  0�      )       P8      B       P                   �      �       0��      �       Q�      �       q�                        "       B        UB       Q        �U�Q       Z        UZ       \        �U�                         "       %        0�(       6        P6       Q        SQ       T        p�T       Z        s�                                     0�               P               p�                      �             U      �       ^�              �U�                      �             T      �       \�              �T�                           �             	��             ]      C       PC      �       ]�      �       P�      �       ]                       �             0�      3       S3      �       1��      �       S�              P                  ,      �       V                      G      N       PN      �       S�      �       U                            \       �        U�       �        S�       �        U�       �        �U��       �       S�      �       �U�                                �       �        P�       �        V�       �        P�       
       V$      7       P7      Z       VZ      _       P_      �       V                      T      e       Ue      �       V�      �       �U�                    T      _       T_      �       �T�                    q      u       Pu      �       S                                   U      S       VS      T       �U�                              #       P#      R       SR      S       v� S      T       �U#h                                �      �       U�      �       �U��      	       U	             \             U              \              �U�             U                    �      �       T�             �T�                        �      �       P�      �       P      =       P             P                  �      �       V                     �             SU      Y       PY      �       S                 �      �       S                      �      �       U�      #       ^#      &       �U�                      �      �       T�      !       ]!      &       �T�                           �      �       	���      �       \�             P             \             P             \                       �      �       0��      �       S�             1�             S      &       P                  �             V                                 P             S                          &      �       U�      �       �U��      �       U�      �       �U��      �       U                          &      �       T�      �       �T��      �       T�      �       �T��      �       T                      &      :       Q:      �       �Q��      �       Q                        -      �       P�      �       P�      �       P�      �       q�                                                    \        U\       g        �U�g       r        Ur       �        �U��       �        U�       �        �U��       K       SK      P       �U�P      �       S�      �       U�      �       �U��      �       S�      �       �U��      �       U                      �       �        P!      #       Pm             P                    }      �       U�      �       �U�                   }      �       9��      �       T                        f      s       Us      x       Sx      |       U|      }       �U�                        �      (       U(      W       SW      ]       �U�]      ^       U                          X       VX      \       r�                    5      8       P8      \       R                    �      �       U�      �       �U�                      R      a       Ua      l       Vl      �       �U�                  �      �       S                   �      �       T�      �       V                   �      �       p A$#���      �       Q                    �      �       P�      �       S                      �      �       U�      M       ]M      R       �U�                  �      F       S                  �      �       \                    �      �       p A$#���      �       Q                    �              P       ?       \                    �      �       U�      �       �U�                    ;      �       U�      �       �U�                 Z      �       P                 l      �       P                              (       U(      5       S5      :       U:      ;       �U�                                      T       6       V6      :       T:      ;       �T�                    
             U             �U�                    
             T             �T�                    �              U       
       �U�                    �             T      
       �T�                        �      �       U�      �       S�      �       U�      �       �U�                        �      �       U�      �       S�      �       U�      �       �U�                        �      �       U�      �       S�      �       U�      �       �U�                                    �       U�      �       �U��      �       U�      �       �U��      �       U�      �       �U��      �       U                    �      K       Pc      i       P                       5       P                      �      �       P�      �       p��      �       P                    N      e       Rm      �       R                                 U             �U�                      �      �       U�      �       �U��      �       U                    �      �       U�      �       �U�                          |      �       U�      �       S�      �       �U��      �       S�      �       U                    �      �       T�      �       T                        @      X       UX      q       Sq      {       U{      |       �U�                 @      N       U                                 2       U2      :       S:      >       U>      ?       �U�?      @       U                      u      �       U�             S      #       �U�                 �             \                  �             V                      �      �       P�             p D@$�      	       P	             R                      �      �       U�      r       \r      u       �U�                        �      �       P�      $       V$      '       P'      p       V                    �      �       P�      t       ]                    �      -       S:      o       S                                   U      R       SR      �       �U�                    I      L       PL      �       V                    .      5       P5      I       V                  _      �       S                      t      ~       U~      �       S�             �U�                    �      �       P�             V                    �      �       P�      �       V                  �             S                        ]      e       Ue      o       So      s       Us      t       �U�                              p      �       U�      J       SJ      S       TS      T       �U�T      V       SV      \       �U�\      ]       U                   �      M       \M      S       U                 �             s8�C%�                                0       U0      j       Sj      n       p�n      o       �U�o      p       U                  J      n       P                        V      s       Us      �       S�      �       U�      �       �U�                    d      �       V�      �       V                  x      �       P                  �      �       \                                     U             S             U             �U�                        �      �       U�             S             U             �U�                    L      U       UU      V       �U�                          �      p       Up              V       )       �U�)      ?       V?      K       UK      L       �U�                 e      p       ^                    i      "       \)      9       \                    m      $       ])      9       ]                    p      �       S)      9       S                   p      &       ^)      9       ^                    |      (       _)      9       _                  �             S                  �      �       S                                    �       U�      �       S�      �       Q�      �       �U��      �       S�      �       �U��      �       U                    �      �       p :#6��      �       �l�:#6�                          ]      o       Uo      y       Sy      }       U}      ~       �U�~             U                        �             U      X       SX      \       �U�\      ]       U                    �      �       P�      W       \                        (       P(      @       p  $1 $+( �                 (      @      ! v �s �DA$"p  $1 $+( �                  k      Y       V                    B      F       PF      k       V                        �      �       U�      �       S�      �       �U��      �       U                  �      �       P                                L      ^       U^      �       S�      �       Q�      �       �U��      �       S�      �       U�      �       �U��      �       U                    u      �       p 8#:��      �       R                          #      5       U5      A       SA      J       UJ      K       �U�K      L       U                                �      �       U�             S             Q             �U�             S      !       U!      "       �U�"      #       U                    �      �       p 6#:�             R                              �      �       U�      �       S�      �       Q�      �       �U��      �       S�      �       �U��      �       U                  �      �       p :#2$�                                      +       U+      e       Se      i       Qi      j       �U�j      z       Sz      ~       U~             �U�      �       U                  J      \       p 8#3�                          �             U             S             U             �U�             U                            �      �       U�      �       S�      �       U�      �       �U��      �       S�      �       �U�                            ^      f       Uf      �       S�      �       U�      �       �U��      �       S�      �       �U�                          �      �       U�      A       SA      \       U\      ]       �U�]      ^       U                    =      I       VI      \       T                  	      M       ]                 =      C       p 5#3�                                    P       K       \K      \       R                        G      x       Ux      �       S�      �       �U��      �       U                     �      �       3 ��      �       4 ��      �       3 �                  �      �       V                  �      �       ]                 �      �       p 5#3�                  �      �       P�      �       ^                          �
      �
       U�
      *       S*      E       UE      F       �U�F      G       U                      �
      &       ]&      2       V2      E       T                 &      ,       p 5#3�                                    P      4       \4      E       R                                        {      �       U�      T	       ST	      X	       UX	      Y	       �U�Y	      �	       S�	      �	       U�	      �	       �U��	      h
       Sh
      o
       Uo
      p
       �U�p
      q
       Sq
      r
       �U�                  �      �       U                            �      �       U�      q       Sq      x       Ux      y       �U�y      z       Sz      {       �U�                      �      �       T�             T             T                    <      >       TN      e       T                      V      �       U�      �       �U��      �       U                    d      �       P�      �       P                   l      �       P�      �       P                 V      ]       U                      >      j       Uj      L       SL      V       �U�                      >      j       Tj      Q       ]Q      V       �T�                       >      j       0�j      �       P�      )       \)      ,       P,      O       \                  j      V       ��                  �             p s8��                         )       P                      �             U      4       S4      >       �U�                            F      �       P�      �       ]�      �       P�             ]      /       P/      9       ]                    I      �       V      /       V                                b      �       �_���      �       �_�^��      �       �8���      &       �^�_�&      =       �^���      �       �^�_��            	 �^�8��            	 �8��_�      /       �8���                  �      �       V                    =      @       P@      >       ��                 =      7       \                      H      ^       U^      b      	 8Hf     b      c       �U�                    H      T       TT      c       �T�                              �        U�       �        �U��       �        U                           �        U�       �        �U�                  6       �        X                  �       �        P                      �       �        U�       A       SA      G       �U�G      H       U                      �       �        T�       B       VB      G       �T�G      H       T                 �       G       0�                   �       B       VB      G       �T�                   �       A       SA      G       �U�                     �       :       ]:      =       }�?      F       ]                  �       ?       \                         9       U                          c      r       Ur      v       �U�v      �       U�      �       S�      �       �U�                 y      �       V                  �      �       P                  �      �       S                      �      �       U�      �       V�      �       �U�                  �      �       V                                    -       p���~�-      8       Q8      ]       S]      g       Qg      �       S�      �       Q�      �       S�      �       ȟ                          �      �       U�      �       �U��      �       U�      �       S�      �       �U�                    �            " u�� $ &2$ [e     "�t u�"�            ( u�� $ &2$ [e     "�u�#<�u�"�                   �            " u�� $ &2$�Ze     "�t u�"�            ( u�� $ &2$�Ze     "�u�#<�u�"�                              %       P%      ^       Vf      �       V�      �       V                  +      �       S                   }      �       0��      �       V                      �      �       U�      �       S�      �       �U�                 �      �       S                        r
      �
       U�
      �
       S�
      �
       �U��
      �
       U                  �
      �
       S                              #      �       U�      �       \�      �       Q�              �U�              \             �U�              U                      #      �       T�             �T�              T                
     #      ,       0�,      w       Q              Q                    *      `       P              P                      o      z       Vz      �       T�             �T�                          l      �       \�      �       Q�              �U�              \             �U�                    �      �       ]              ]                    �      �       ~ p "��      �       T                   �      �      	 | �#�� ��      �       Q                          �      �       P�      �       S�      �       U              S             U                        z      �       V�              �TC%�              V             �TC%�                  �      �       S                          ^      w       Uw      `       V`      d       Ud      e       �U�e      f       U                        n      w       Uw      `       V`      d       Ud      e       �U�                    1      5       P5      _       S                  �      �       P                    �      �       P�      1       S                  �      %       P                        %       R                      �             U      �       w �      �       ��                      �             T      �       ]�      �       �T�                               �             	��      "       V"      O       PO      "       V"      &      	 r z ��&      w       ������w             V      �       P�      �       V                    �      &       Y&      o       ��o             Y                     �      �       0��             Qw      z       q�                     �      �      
 r8z ���      �       q 3$s� "#8z ���      &      	 r z ��&      w       ������                 �      �      	 { 0$0&�                   �      o       0�o      w       1�w             0�                       �             0�      ?       ^?             1�      �       ^�      �       P                      8      "       S"      &       R&      o       ��o      w       Rw             S                     �      �       r8�      &       R&      w       ��                          S      Z       PZ      �       ^-      1       P1      r       Sr      w       r�                      �             0�      �       \�      �       \                       �             0�      �       _�      �       _�      �       _                      �      �       U�      �       w �      �       ��                      �      �       T�      �       \�      �       �T�                           �      �       	���      �       S�             P      �       S�      �       P�      �       S                       �      �       0��      �       V�      �       1��      �       V�      �       P                  �      G       Vr      �       V                        �             X      �       ]�      �       P�      �       ]                                 P      �       ^                 �      �       �����      >       _                    �      �       P             P                              <        U<              S      	       �U�                                        8        T8       G        �T�G       M        TM       �        �T��       �        T�       �        �T��       �        T�       	       �T�                                                <        Q<       G        �Q�G       \        Q\       j        �Q�j       r        Qr       �        �Q��       �        Q�       �        �Q��       �        Q�       �        �Q��              Q      	       �Q�                                                  <        R<       G        VG       \        R\       j        Vj       r        Rr       �        V�       �        R�       �        V�       �        R�       �        V�              R             V      	       �R�                                              X       <        X<       G        �X�G       \        X\       j        �X�j       r        Xr       �        �X�                                    !        Y(       <        Y<       G        �Y��       �        Y�       �        Y�       �        �Y�                          =       ?        P]       _        Ps       u        P�       �        P�       �        P                     4       G        \Q       j        \j       �        \�       �        \�              \                          	      #       U#      �       S�      �       �U��      �       S�      �       �U�                      *      7       P7      �       V�      �       V                    J      �       S�      �       �U�                                          �       U�      ;       S;      H       TH      I       �U�I      �       S�      �       U�      �       �U��      	       S	             �U�             U                                    �       T�      �       X�      3       ��3      �       �T��             T             �T�             T                                          �       Q�      @       ]@      H       UH      I       �Q�I      �       ]�      �       u��      �       �Q��             Q             �Q�             Q                                 u       Ru      �       V�      <       VI      �       V�             R             R                    �      �       P�      3       ^                   �      �       P�      �       Q�      �       P                      a      >       \I      �       \�             \                    �      �       P�      3       _                 �             v  $d $-( �                    \	      3
       U3
             �U�                      \	      �	       T�	             S             �T�                  �
             R                               P                                                                                                                    
      T       UT      s       \s      �       U�      �       \�      #       U#      @       \@      H       UH      {       \{      �       U�      �       \�      4       U4      >       \>      S       US      p       \p      z       Uz      �       \�      �       U�      �       \�      �       U�      �       \�      �       U�             \      "       U"      ?       \?      L       UL      i       \i      v       Uv      �       \�      �       U�      �       \�      �       U�             \             U      3       \3      =       U=      Z       \Z      d       Ud      ~       \~      �       U�      �       \�      �       U�      �       \�      �       U�      �       \�      	       U	      Q	       \Q	      V	       �U�V	      Z	       \Z	      [	       �U�[	      \	       U                                                                                                                                  
      Q       TQ      s       �T�s      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�              �T�              T             �T�              T       @       �T�@      E       TE      {       �T�{      �       T�      �       �T��      4       T4      >       �T�>      P       TP      p       �T�p      r       Tr      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�             �T�             T      ?       �T�?      I       TI      i       �T�i      s       Ts      �       �T��      �       T�      �       �T��      �       T�             �T�             T      3       �T�3      :       T:      Z       �T�Z      a       Ta      ~       �T�~      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      
	       T
	      [	       �T�[	      \	       T                 $      3       t�                        �      �       V�      �       T�      �       v��      �       V                          ;       P[	      \	       P                                                   $      0        �0      5       ]�5      n        �n      s       ]�s      �        ��      �       ]��      �        ��      �       ]��              �             ]�               �       "       ]�"      4        �4      >       ]�>      �        ��             !�      .        �.      3       !�3      U        �U      Z       !�Z      |        �|      ~       !�~      �        ��      �       !��      �        ��      �       !��      �        ��      �       !��      	        �	      O	       VO	      U	       T                U      w       1�                U      w       d�                |      �       2�                |      �       ȟ                {      �       0�                �      �       1�                �      �       1�                �      �       2�                �      �       3�                             4�                "      )       5�                    5      F       TF      ^       �T�                      1      l       Ul      /       S/      5       �U�                                1      l       Tl      t       ]t      �       T�      �       ]�      �       T�      *       V*      4       ]4      5       �T�                            1      `       Q`      �       �Q��      �       Q�      �       �Q��      �       Q�      5       �Q�                  �      &       P                         !       1�!      *       Q                                        U       *       S*      .       �U�.      1       U                                %        T%       +       V+      .       �T�.      1       T                                    %        Q%       S        \S       U        PU       _        \_       o        P.      1       Q                 m       )       T                  �       )       \                  �       )       V                  �       )       S                  a      t       Q                        �      �       T�      �       �T��             T      
       �T�                 �      �       1�                 �      �       U                      O      `       U`      �       V�      �       �U�                    i      p       Pp      �       S                    �      �       U�      N       ^N      O       �U�                  �      �       T�      H       V                 �      L       ]                          4       \4      7       |�                  �      G       S                  &      /       P                       %      	 | 3$s� "                    q      �       U�      �       ^�      �       �U�                       �      �       0��      �       \�      �       |��      �       \                 �      �       ]                  �      �       V                  �      �       S                  �      �       P                 �      �      	 | 3$s� "                      1      :       U:      p       Vp      q       �U�                           1      :       	��:      F       SF      j       Pj      m       Sm      n       Pn      o       S                  X      j       U                      �      �       U�      ,       V,      1       �U�                      �      �       T�      0       ]0      1       �T�                      �      �       Q�      .       \.      1       �Q�                    �      �       P�      +       S                      C      [       U[      �       V�      �       �U�                    f      j       Pj      �       S                      �              U      B       VB      C       �U�                                 P      A       S                         *        U                  8       X        U                        x       �        U�       �        S�       �        �U��       �        U                      �       �        U�       �        S�       �        �U�                  �       �        Q                        �       �        U�       �        S�       �        �U��       �        U                      �       �        U�       �        S�       �        �U�                            /       U/      ^       V^      a       �U�                          /       T/      a       �T�                  /      W       S                        8      K       \K      O       TO      P       |�P      V       \                  �      �       U�             �U�                  �      �       T�             �T�                  �      �       Q�             �Q�                        �             ^             U             ~�             ^                 �             S                  �             V                  �             ]                 �      �       S                  �             \                  �      �       R�             �Q@$�                    E      Z       UZ      �       �U�                  g      �       P                 g      �       U                 g      �       T                        �      �       U�      5       Y5      D      	 XJf     D      E       �U�                        �      �       T�      �       T�             X      E       �TC%�                      �      &       Q&      D      	 PJf     D      E       �Q�                      �      )       R)      D      	 tIf     D      E       �R�                      �      �       X�      D      	 �Jf     D      E       �X�                        D       [                        D       Z                      %      3       U3      4       �U�4      �       P                        %      3       T3      4       �T�4      Z       SZ      �       X�      �       �TC%�                      %      3       Q3      �       V�      �       �Q�                  �      �       Q                  �      �       R                                �             U             V      �       �U��      >       V>      j       �U�j      �       U�      �       V�      �       �U�                        O      S       | p "�S      �       | ~ "�>      b       | ~ "�      �       ^                        _      c       } p "�c      �       }  "�>      b       }  "�       �       _                            }      �       P�      �       Q>      a       Q:      >       P>      Q       QT      d       Q                      6      �       V>      b       V�      �       ]                   �      �       S�      b       S                   j      �       u�      �       v                      �      �       P             P0      >       P                          �      �       P�      �       \�      >       \�      �       P�      �       ]                  �      �       P                  �      �       P                                  t      �       U�      �       \�      �       U�      B       \B      K       UK      R       �U�R      c       Uc      �       \�      �       �U�                 �      B       S                     B      K       uR      c       uc      g       |                    �      �       P      +       P                    �      �       P�      �       \�      �       q  $|  $-( �                 �      �       P                       �      �       P�      -       Vy      }       P}      �       ]                          7      [       U[      �       S�      �       U�      �       �U��             S      %       �U�                  �             \                      �      �       T�      g       V�      �       V                    �      �       Z�             ��                  �             _                    �      �       P�      �       V                  �      �       P                     [      [       3} �[      ^       4} �^      `       3} ��             4} �                      �      �       U�      s       Vs      t       �U�                  �      r       S                      (      @       U@      v       Sv      �       �U�                  <      z       |  $v  $)��                                        �        U�       �        �h�       g       Ug      �       �h�      �       U�      �       �U��      �       U�      �       �U�                            9       �        R�       �        R�       !       t� �u� �"�!      g       @Jf     #h�u� �"��      �       R�      �       R                    �       �        p 8#t�#L��y      |       p 8#t�#L��                      �	       
       U 
      ,       ^,      /       �U�                        �	      
       T
      +
       U+
      .       _.      /       �T�                          �	      �	       Q�	      

       R

      
       Q
      +
      	 xIf     +
      /       ��                 �
      �
       S                  �
      &       V                  �
      (       \                  �
      *       ]                 �
      %       S                      �
      �
       X�
      �
       ���
      �
       X                  ,
      F
       P                      �             U      	       �U�	             U                      �             U      	       �U�	             U                    �      �       R	             R                              X       UX      a       Sa      �       �U��      �       U                    r      a       Sa      �       �U�                         a       Sa      �       �U�                  w      �       S                    2      M       PP      Z       P                          �      �       U�      �       �U��      	       U	      (	       S(	      ,	       �U�                   	      	       0�	       	       p  $@L$)��                 �      �       �U�                        ,	      �	       U�	      �	       V�	      �	       �U��	      �	       U                      G	      �	       U�	      �	       V�	      �	       �U�                  Q	      �	       u�t��                 Q	      �	       u�t��                     Q	      s	      $ u�t� $u�t� $+( �s	      {	       s @&�{	      �	       S                      /      W       UW      �      	 @Jf     �      �       �U�                      /      Z       TZ      �       P�      �       �T�                    /      �       Q�      �       �Q�                  �      �       P                  �      �       �U�                  �      �       �T�                  �      �       �Q�                        "       S|      �       S                            A       VE      p       V�      �       \                    "      "       P"      h       ]�      �       ]                     "      A       \E      a       \�      �       V                  "      Z       S�      �       S                    )      N       ^�      �       ^                      �      �       U�             S      (       �U�                      �      �       T�      �       V�      (       �T�                            �      �       Q�      &       ^&      6       s6      L       �Q�L      �       ^�      (       �Q�                          �      &       ^&      6       s6      L       �Q�L      �       ^�             �Q�                    �      �       V�             �T�                  �             S                          L       \�             \                          L       ]�             ]                      �      �       P�      �       _�             _                    �      �       P�             P                    �      �       V�             V                      �      �       U�      .       S.      X       �U�                    �      .       S.      O       �U�                    '      +       P+      O       V                      X      �       U�      �       S�      7       �U�                    �      �       S�      7       �U�                    �      �       P�      �       \                    �      �       P�      .       V                  �      �       P                    �      �       P�      �       S                  �             P                                 P      6       \                     �      L       UL             U      �      	 �Vf                           �      g       Tg      �       T�      �      	 �Vf     �      4	       V                     �      o       Qo      t       ^t      �       �Q�                     �      q       Rq      v       Sv      �       �R�                    �      &       X&      `
       ��                    �      U       YU      `
       ��                            �      �       T�      �       ���      �       T�      	       ��	      *	       T*	      �	       ��                 �      �	       ]                           �      �       Q�      �       ���      	       Q	      	       ��	      *	       Q*	      `
       ��                            �      �       R�      �       ���      	       R	      	       ��	      *	       R*	      `
       ��                        j	      l	       P�	      �	       P�	      A
       SO
      V
       S                      �      �       P	      	       P*	      `
       ��                              �      �       _�      	       _*	      >	       _X	      l	       Vv	      �	       V�	      �	       V�	      �	       U                    �	      D
       \O
      Y
       \                    >	      J
       _O
      _
       _                   �	      
       ��
      `
       ��                   �	      F
       ]O
      [
       ]                    �      �       1��      	       	��*	      `
       ��                      E	      l	       1�n	      �	       	���	      H
       ^O
      ]
       ^                         �	      �	       0��	      .
       @v �.
      0
       Av �0
      2
       @v �O
      W
       @v �                                        U       <        P<       n        �U�n       t        P                              X        TX       ^        �T�^       t        T                                       0�               U       &        Qn       s        Q                                         0�       H        X^       d        Xn       q        Xs       t        X                      B       L        p 2�L       Q        P^       h        p 4�h       n        P                  4       n        R                      �      �       U�      �       ]�      �       �U�                      �      �       T�      �       V�      �       �T�                       �      �       �Jf      Kf     @��      �       s��      �       S�      �       s�                  �      �       Q                  �      �       P                     �      �       0��      �       \�      �       \                      $      s       Us              ]              �U�                  h             ^                  h      �       \                  h             ��                  h      �       S                    �      �       P�             _                  �      �       P                 $      w        �Vf     ��Vf     �' $0+��                  �      �       P                 �      �       T                 �      �       U                            T       UT      "       S"      $       �U�                        `      d       Pd      p       V�      �       P�      #       V                    n      p       P�      �       P                  �             P                              T                              U                      4      f       Uf      �       �U��      �       U                      4      f       Tf      �       �T��      �       T                        4      ^       Q^      �       V�      �       �Q��      �       Q                  f      �       S                      �      �       U�      .       �U�.      4       U                      �      �       T�      .       �T�.      4       T                        �      �       Q�      -       V-      .       �Q�.      4       Q                  �      ,       S                                 U!      %       U                      �      	       U	      �       S�      �       �U�                            ,       P,      �       s� �      �       �U#X                         =       R                        K      N       p G&�N      U       PU      �       Q�      �       Q                  �      �       Q                      �      �       p G&��      �       P�      �       Q                          -       Q-      ^       u8                          $       R$      ^       u�                           �      �       U�             ]             �U�             ]             �U�                          �      �       T�             S             �T�             S             �T�                    �             | p "�             U                        �      �       v p ��             V             T             V                            ^       U^      �       �U��      �       U                            B       TB      �       �T��      �       T                              j       Qj      �       S�      �       �Q��      �       Q                  ?      [       R                    K      c       Tc      �       V                    v      }       P}      �       \                  ~      �       P                    5      �       U�      �       S�             �U�                        5      �       T�      �       \�      �       T�      �       \�             �T�                                           5      q       0�q      �       r  $p  $+���      �       r  $t #� $+���      �       r  $p  $+���      �       v ���      �       0��      �       r  $p  $-���      �       r  $p  $-���      �       v ���      �       0��      �       P�      �       0��      �       P�              V                                 5      q       0�q      �       p  $q  $-���      �       t #� $q  $-���      �       p  $q  $-���      �       t #� $q  $-���      �       0��      �       p  $q  $+���      �       p  $q  $+���      �       t � $q  $+���      �       0��      �       P                          �       �        U�       �        �U��       �        U�       �        �UO&�U'�UO&��       �        U                        �       �        T�       �        �T��       �        T�       �        �TO&�T'�TO&�                      t       z        Uz       �        u���       �        �U�                    t               T       �        Z                  �       �        Y                      �              U      4       �U�4      5       U                      �              T      4       �T�4      5       T                        �              Q      '       S'      4       �Q�4      5       Q                                T      (       V                    !      %       P%      -       \                  &      0       P                    �       �        T4      5       T                    �       �        Q4      5       Q                    �       �        U4      5       U                      -      K       UK      9       \9      B       �U�                      -      E       TE      =       ^=      B       �T�                      �      �       P�      7       V7      A       U                      C      _       V_      �       S�              v8                 �      �       |                 �      �       |                   �      �      	 | �@A$"��      �       Q                            W      m       Pm      y       ]y      �       P�      �       ]�      �       P�      �       0��      ;       ]                      '      @       U@      &       V&      -       �U�                      '      =       T=      *       ]*      -       �T�                      '      G       QG      K       RK      -       �Q�                      O      V       PV      %       S%      -       P                    �      �       P�      (       \                      �             P
      
       P
             p  $1 $+( �             r  $1 $+( �                  �      &       U&      '       P                            �      �       U�      �       S�      �       U�      �       �U��      �       S�      �       �U�                                 U      �       �\                                   T      L       w L      �       �T�                                     Q      '       \'      5       s p :$| "�<      @       Q                                         R      �       V�      �       p	��      �       �R��      �       V�      �       p	�                          A      P       PP      �       w �      �       �P�      �       w �      �       �P                          �       U�             �\                          �       T�             �X                              �       Q�      �       V�      �       s p :$v "��      �       Q                        �      �       P�      �       S�      �       U              S                            �
             U             �U�      Z       UZ      |       S|      ~       �U�~             U                      `      h       Ph      k       p�k      w       r�                    C      E       PJ      U       P                                 P      z       V                  �      �       U                  �      �       T                  �      �       Q                        V	      �	       U�	      �
       V�
      �
       �U��
      �
       U                  �	      �
       \                   �	      �	       v �0$0&@$��	      �	       U                   �	      �	       v�0$0&@$��	      �	       T                 �	      �
       @K$�                    �	      �	       P�	      L
       R                            V
      ]
       0�]
      d
       1�d
      k
       2�k
      r
       3�r
      y
       4�y
      �
       5�                  �      M	       V                  �      M	       \                  �      	       Q                  �      �       P                      �      �       P	      -	       P-	      M	       R                 c      �        Wf     � $ &: Yf     "�                       �      �       0��      �       P�      �       p��      �       r�                        +      �       U�      �       S�      �       U�      �       �U�                              
        U
       *       ^*      +       �U�                                      T       (       ](      +       �T�                                      Q       $       V$      +       �Q�                              #        R#       &       \&      +       �R�                      ,       .        P.       #       S#      +       P                                  l      �       U�      �       S�      �       U�      �       �U��             S      !       U!      "       �U�"      #       S#      $       �U�                            [      �       U�      _       S_      f       Uf      g       �U�g      h       Sh      l       �U�                    t      `       Vg      i       V                    x      b       \g      k       \                               Q                  �      �       P                        �      �       P�      �       P             P      f       R                     �      _       s��_      f       u��f      g       �U#��                            �      �       U�      �       S�      �       U�      �       �U��      $       S$      &       �U�                  
      A       P                                           q r �      #       Q#      )       s� �1&r t �"�)      /       s� �1&s �t �"�/      4       Q4      >       s� �1&r t �"�>      A       s� �1&s �t �"�                  O      �       v ����5+��                            3      Z       UZ      �       S�      �       U�      �       �U��      �       S�      �       �U�                      �      �       U�      1       S1      3       �U�                        �      �       T�             T      (       V(      /       T                    �             P             s�                                  &      ]       U]      ^       �U�^      �       U�      I       SI      T       UT      U       �U�U      R       SR      Z       �U�Z      [       U                            ^      �       U�      I       SI      T       UT      U       �U�U      R       SR      Z       �U�                    �      �       T�             T                    �      �       Q�             Q                    p      N       ]U      W       ]                        �      �       \�      �       P�      �       \�      �       0��      L       \U      U       \                        �      �       V�      �       P�      �       V�      �       0��      J       VU      S       V                        �      �       U�      �       �U��      �       U�      �       �U�                         �      �       0��      �       P�      �       S�      �       p��      �       s�                    n       �        U�       �        �U�                     n       p        0�p       �        P�       �        p�                     2       4        0�4       d        Qd       g        q�                                   0�       (        Q(       +        q�                      �       �        U�       x       Vx      �       �U�                      �       �        T�       ~       ^~      �       �T�                      �       �        Q�       �        _�       �       �Q�                                   P      f       Sf      j       U                           �       �        	���       �        ]�              P      p       ]p      v       Pv      |       ]                       �       �        0��       �        S�       p       1�p      w       Sw      �       P                    �              R      p       _                                �              U       �       S�      �       U�      �       �U��      �       S�      �       �U��      �       S�      �       �U�                            
       P
      �       V�      �       P                      N      V       UV      �       S�      �       �U�                     U      V       0�V      �       V�      �       v�                      U      V       u��V      �       v Hs "#���      �       v Hs "#��                  b      �       R                    *      M       UM      N       �U�                     *      5       0�5      C       1�C      N       2�                                  U       *       �U�                          %       T%      *       �T�                      �
      �
       U�
             V             �U�                 �
      �
       0�                     �
      �
       ?} ��
      �
       @} ��
             ?} �                 �
      �
       0��
             \                   �
      �
       v8�s "@I$��
      �
       T                          �	      �	       U�	      X
       SX
      ^
       �U�^
      `
       S`
      b
       �U�                          �	      �	       T�	      Y
       VY
      ^
       �T�^
      a
       Va
      b
       �T�                      �      �       U�      �	       S�	      �	       �U�                    �      �       T�      �	       �T�                     >	      �	       D~ ��	      �	       E~ ��	      �	       D~ �                    M	      f	       \f	      �	       V                    F	      I	       p 3#5�I	      �	        3#5�                      a      t       Ut      �       S�      �       �U�                    a      g       Tg      �       �T�                     �      �       7v ��      �       8v ��      �       7v �                      �      �       U�      \       S\      a       �U�                    �              T       a       �T�                        �      �       U�      �       \�      �       U�      �       �U�                      �      �       T�      �       S�      �       �T�                   �      �       V�      �       T                    �      �       X�      �       �\                      *      >       U>      �       V�      �       �U�                          3      O       SO      U       s��� �U      a       Ta      r       s��� �r      x       s���`�x      �       T�      �       s���`�                      �             U      $       S$      *       �U�                    �      �       T�      *       �T�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                          �      �       U�             V             �U�      �       V�      �       �U�                    �      �       T�      �       �T�                              �      �       ]�             S      :       S:      X       PX      a       p���g�c      n       Pn      w       p���                      �      �       p :#1$��      	       | :#1$�      �       | :#1$�                    �      �       P�      �       R                      �      �       U�      �       V�      �       �U�                    �      �       T�      �       �T�                          3       \3      m       S                                 X      �       �\                  :      P       P                        �      �       U�      �       S�      �       U�      �       �U�                    �      �       T�      �       �T�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                          J      x       Ux      y       �U�y      �       U�      �       �U��      �       U                          J      t       Tt      y       �T�y      �       T�      �       �T��      �       T                    E      I       UI      J       �U�                    E      I       TI      J       �T�                              5       U5      6       �U�6      D       UD      E       �U�                              5       T5      6       �T�6      D       TD      E       �T�                                        #       U#      y       Sy      �       U�      �       �U��      �       S�      �       U�      �       �U��             S             �U�                                    ?       T?      |       \|      �       �T��      �       \�      �       �T��             \             �T�                    �      �       v 
���      �       q 
��                                 U             �U�                        	      +       U+      _       S_      c       Uc      d       �U�                  J      c       Q                    �       �        U�       	       �U�                 �       �        u(                             $        U$       �        V�       �        �U�                             $        T$       ,        ],       �        �T�                           {        Q�       �        Q                    $       �        \�       �        �T $ &H�U"#��                      K       e        Pe       �        r��       �        r�                      d      �       U�      �       �U��      �       U                    q      �       T�      �       T                   �      �       R�      �       R                          �      �       U�      �       S�              �U�              S             �U�                    �      �       S�              �U�                                                 P�      �       P3      7       P�      �       Pk      o       P�      �       P@      D       P�      �       P�      �       T�      �       P                    0      4       P4      �       S                    �      �       P�      3       S                    O      S       PS      �       S                    �      �       P�      k       S                    �      �       P�      �       S                    �      �       P�      @       S                   \      `       P`      �       S                   0      4       P4      �       S                  B      H       P                   �      �       P�             S                  �      �       P                   O      S       PS      �       S                  i      o       P                   �      �       P�      D       S                  �      �       P                   �      �       P�      �       S                  �      �       P                   �      �       P�      >       S                  �             P                   \      `       P`      �       S                  f      l       P                    �      �       S�      �       S                    �      �       P�      �       p�                 �      3       S                 J      �       S                 �      "       S                 F      �       S                 �      �       S                        @      T       P�      �       P�      �       T�      �       P                            )       U,      0       U6      :       U                        6       S                    l      p       Pp      �       S                   l      p       Pp      &       S                      �      �       P�      �       p��      �       P                 �      !       s��                  (              S                 R      �       S                 r      y       s(                 z      �       s0                 �      �       s�                  �      �       s�                  �      �       s�                  �             s�                 Z      d       s�                 �      �       s��                 �      �       s�                                    0�      *       V*      t       v�t      ~       V~      �       0��             \                            .       S.      |       s��|      �       S                  �             V                  �      �       S                         
      *
       0�*
      6
       V6
      x
       v�x
      z
       Vz
      �
       0��
             \                      *
      :
       S:
      x
       s��x
      �
       S                  �
             V                  �
      �
       S                 ]      l       0�                                        '      3       V3      6       v�>      J       VJ      M       v�`      l       Vl      o       v��      �       V�      �       v��      �       V�      �       v��      �       V�      �       v�}	      �	       2} ��	      �	       3} �                  �	      �	       P                 �      �       0�                            �      �       V�      �       V�      �       V�      �       V             V      )       V�      $       2} �$      '       3} �                  �      �       p ��                            �      �       0��      �       Hs ��      �       Is ��      �       Hs ��      �       s w @�J      Y       SY      \       s�                  j      r       S                  u      }       V                 z      �       P                      �      �       U�      �       \�      �       �U�                               �      �       0��      �       S�             V             S             V             v�             V=      C       s w �s      ~       S                      �       �        U�              S      	       �U�                      �       �        U�       �        S�       �        �U�                 �       �        u                  �       �        s                   �       �        s��       �        �U#�                   �       �        s�       �        U                      �             U      "       S"      #       �U�                         "       s�"      #       �U#�                       !       P                  !      2       S                     !      )       V)      .       v�.      3       V                 �      �       P                  �      �       S                 �      �       V                        d       k        Uk       }        S}       �        U�       �        �U�                     �      �       \�      �       v �8$| !��      �       V                    R       Y        UY       d        �U�                      �      �       S�      �       p �8$s !��      �       P                      [      s       Us      �       S�      �       �U�                                    U       #        u                         .
      �
       U�
      �
       S�
             sP�      �       �U�                    .
      �
       T�
      �       ��                    .
      �
       Q�
      �       �Q�                    .
      7
       R7
      �       �R�                    �      �       S�      �       s�                      /      6       P6      �       V�      �       |w�                 x      o       \                    �      �       S�      �       U                 �      �       ]                  �      o       S                    �      c       ]c      o       }p�                       �      	       0�	             Q             R      %       q�%      A       Q                       	             q 3�             r 3�             R      A       q3�                     �      	       ]	             P      %       p�%      C       P                    h      m       p��m      o       p��                  �      �       P                                                0�      H       QH      O       0�O      �       T�      �       0��      �       R�      �       r��      �       R�      '	       T'	      *	       t�,	      .	       T.	      )
       V                   E	      Y	       \z	      #
       \                      H      �       Q�      ,	       PV	      z	       ]                        �      	       R	      '	       Q.	      
       S
      
       s��
      (
       S                                   P      /       pp�/      ?       P                                p
�0$0&8u "�      /       pz�0$0&8u "�                            �	      �	       P�	      �	       s �	      �	       t G&��	      �	       t G& $0 $+( ��	      	
       P	
      
       s,
      
       r G&�
      
       r G& $0 $+( �                      Z      a       Ua      �       S�      �       �U�                   b      o       p 2��      �       S                  b      o       P                        x      �       U�      Q       VQ      Y       UY      Z       �U�                  �      �       P                     �      �       0��      �       ]�      5       }�5      U       ]                      �      �       P�      $       s|�$      5       s^�L      P       s|�                      �      �       \�      J       |h�J      S       \                        �      �       U�      m       \m      w       Uw      x       �U�                 O      O       P                 O      o       ]                 O      O       PO      k       V                 O      j       S                  �      e       _                  �      e       ^                      <      T       UT      �       V�      �       �U�                   Z      ^       P^      n       S                     n      �       \�      �       |��      �       \                     n      �       S�      �       sv��      �       S                  n      n       Pn      �       ]                 s      �       1�                        q      x       Ux      7       S7      ;       U;      <       �U�                  �      �       P                   �      �       0��      ;       T                     �             0�      (       1�(      4       2�                  �      �       0�             0�                 �      ;       P                  �      ;       Q                        �      �       U�      j       \j      p       Up      q       �U�                  �      �       P                     �      �       0��             ]      `       }�`      l       ]                      �      �       P�      3       s|�3      `       sb�b      g       s|�                    �             V      `       v��`      h       V                        
             U      �       S�      �       U�      �       �U�                    T      V       PV      �       T                     e      k       0�k      v       Qv      |       q�|      �       Q                       T      V       PV      k       Tk      |       t p "�|      �       t p "#��      �       t p "�                        e      k       Rk      |       p 2$r "�|      �      
 p 2$r "#��      �      
 p|2$r "#��      �       p 2$r "�                        �       �        U�              V      	       U	      
       �U�                 +      +       P                 +             ]                 +      +       P+             \                 +              S                        �      �       P�      �       P�      �       s �      �       P                 �      �       |�0$0&�                    �      �       Q�      �       Q                                        U       k        Sk       o        Uo       p        �U�                  :       o        P                       A       I        0�I       c        Qc       f        q�h       o        Q                         :       I        PI       c        q 2$p "�c       f       
 q 2$p "#�f       h       
 q2$p "#�h       o        q 2$p "�                          A       I        TI       c        q 3$t "�c       f       
 q 3$t "#�f       h       
 q3$t "#�h       o        q 3$t "�                      U             U             �U�      #       U                      U             T             �T�      #       T                    `      i      
 p r ��i      �       u� r ��                 `      �       t� r ��                    �      �       P�      �       Q                     �      �       p 3&��      �       q 3&��      �       Q                   �      �       1p 7$��      �       1q 7$�                           �      �       U�      �       �U��      �       U�      �       �U��      �       U�      U       �U�                      �      $       S$      Q       QQ      S       S                        �      �       P�      '       V'      G       v 1'�L      T       V                      �       �        U�              S      �       �U�                  $      �       S                      1      =       YF      �       Y�      .       Y                          u             P      �       ]�      �       P�      �       Z�      .       Z                      �      �       P�      �       P�      �       P                        �       ^                               S                  �      �       \                 �      �       _                        �       V                        �       ]                  M      e       P                  V      r       [                      1      4       P4      M       QM      `       ��                    N      `       Pz      �       P                          h       |        U|       �        ]�       �        �U��       �        ]�       �        �U�                          h       y        Ty       �        S�       �        �T��       �        S�       �        �T�                    �       �        | p "��       �        U                        �       �        v p ��       �        V�       �        T�       �        V                            G        UG       h        �U�                            J        TJ       h        �T�                     B       G        u q ��G       P        UP       g       	 �Uq ��                   B       J        t x �J       g        �Tx �                  V       g        U                  [       g        T                                 T                                 Q                                 U                  �      e       S                               �      �       0��      c       Vc      e       0�e      �       S�      �       s��      �       S�      �       P�      �       p��      �       P�      �       p�                    B	      \	       U\	      f       ��                  �	      T       S                        �	      �	       P�	      �	       ^�	      �	       P�	      T       ^                      �	      �	       Q�	      �	       Q�
      �
       Q                       B	      \	       	��\	      l	       \l	      �	       P�	      _       \                   B	      \	       0�\	      �	       Z�	      T       1�                    �	      �	       P�	      �	       P                       �
      �
       P�
             V             P      I       V                   �
      �
       _�
      I       _                   �
      �
      	 ��e     �
      I       ]                 �	      �
       ��                 �	      �
       S                 �	      �
       �*�	                   �	      �
       ��	                      4
      I
       PI
      Y
       p�                        i       R                  A      U       Q                                         r       P       TP      S       t�U      [       Tk      �       P�      �       p��      �       P                      w      �       Q�      �       p 3$�cf     "�      �       p3$�cf     "                                  	             U      n       Sn      s       �U�s      �       S�      �       �U��      �       S�      �       �U��      �       S�      �       �U�                                    k       Qk      m       u� s      y       Q�      �       Q�      �       Q�      �       u� �      �       Q                              �      �       U�      �       �U��      �       U�      �       �U��      �       U�             �U�      	       U                            �      �       T�             S             U             �T�             S      	       T                 �      �       0�                    X      �       U�      �       �U�                                                                                                                                                                                                                                                                                                    X      �       T�      �       �T��      �       T�             �T�             T             �T�             T             �T�             T             �T�             T      !       �T�!      (       T(      -       �T�-      /       T/      1       �T�1      6       T6      8       �T�8      =       T=      ?       �T�?      F       TF      L       �T�L      N       TN      S       �T�S      Z       TZ      _       �T�_      d       Td      i       �T�i      n       Tn      s       �T�s      x       Tx      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�             �T�             T             �T�             T             �T�             T      %       �T�%      *       T*      /       �T�/      4       T4      6       �T�6      =       T=      G       �T�G      L       TL      M       �T�M      ]       T]      `       �T�`      e       Te      o       �T�o      t       Tt      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T��              T              �T�      	       T	             �T�             T             �T�             T             �T�             T             �T�      $       T$      &       �T�&      +       T+      -       �T�-      2       T2      4       �T�4      ;       T;      =       �T�=      B       TB      D       �T�D      I       TI      K       �T�K      P       TP      U       �T�U      Z       TZ      _       �T�_      d       Td      i       �T�i      p       Tp      y       �T�y      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T�                                                                                                                                X      �       Q�             �Q�      #       Q#      -       �Q�-      F       QF      L       �Q�L      U       QU      _       �Q�_             Q      �       �Q��      �       Q�      �       �Q��      �       Q�      �       �Q��      �       Q�      �       �Q��      �       Q�      �       �Q��      �       Q�      �       �Q��      �       Q�             �Q�      "       Q"      %       �Q�%      8       Q8      G       �Q�G      L       QL      M       �Q�M      ]       Q]      `       �Q�`      e       Qe      o       �Q�o      {       Q{      �       �Q��      �       Q�      �       �Q��      �       Q�      �       �Q��      �       Q�      �       �Q��      �       Q�      �       �Q��      �       Q�             �Q�             Q             �Q�             Q             �Q�      6       Q6      =       �Q�=      k       Qk      y       �Q�y      �       Q�      �       �Q��      �       Q�      �       �Q�                                                      n      �       S�      H       SM      �       S�      �       U�      �       S�      �       U�      �       S�      �       U�      �       S�      �       U�             S             U      t       St      x       Uy      �       S�      �       U�      �       S�      �       U�      �       S                 �      �       0�                        "      -       U-      G       XG      U       TU      X       X                    "      -       T-      X       �T�                       "      -       0�-      P       RP      S       r�U      X       R                   "      -       T-      X       Q                 2      A      	 r 3$x� "                  B      K       P                      �      �       T�              t�       "       �T�                     �      �       t��              T      !       P                        �      �       U�      �       X�      �       T�      �       X                       �      �       0��      �       R�      �       r��      �       R                 �      �      	 r 3$x� "                  �      �       P                   �      �       0��      �       Q                        �      �       U�      �       X�      �       T�      �       X                       �      �       0��      �       R�      �       r��      �       R                 �      �      	 r 3$x� "                  �      �       P                   �      �       �����      �       Q                              �             U      !       ]!      =       T=      @       ]@      C       TC      |       ]|      �       �U�                      �             T      \       V\      �       �T�                	           �             0�      O       \O      R       |�T      \       \\      ^       1�^      a       p�n      p       p�                	     �             0�      C       SC      K       s�K      w       S                  \      p       V                 	            	 | 3$}� "                          #       P#      T       ^                   �             T      �       _                        �      �       U�      �       X�      �       T�      �       X                       �      �       0��      �       R�      �       r��      �       R                 �      �      	 r 3$x� "                  �      �       P                   �      �       ���p��      �       Q                        }      �       U�      �       X�      �       T�      �       X                             �       0��      �       R�      �       r��      �       R                 �      �      	 r 3$x� "                  �      �       P                        �       Q                    F      P       UP      g       �U�                          !       U!      F       �U�                    �       �        U�              �U�                      &       b        Vb       f        Uf       �        V                  *       �        \                                                                                                                        k      �       U�      �       Q�      �       �U��      �       Q�      �       �U��             Q             �U�             Q             �U�      !       Q!      #       U#      (       Q(      0       U0      7       �U�7      @       Q@      G       UG      I       QI      P       UP      \       Q\      _       �U�_      z       Qz      �       �U��      �       Q�      �       �U��      �       Q�      �       �U��      �       Q�      �       U�              Q              �U�             Q      *       �U�*      3       Q3      6       �U�6      S       QS      Z       UZ      j       Qj      l       Ul      q       Qq      x       Ux      �       Q�      �       U�      �       Q�      �       U�      �       �U��      �       Q�      �       �U��      �       Q�      �       �U��      �       Q�             �U�             U                        k      �       T�             S             �T�             T                    k      �       Q�             �Q�                                  @       U@      _       V_      e       Ue      f       �U�f      h       Vh      k       �U�                                ,       T,      a       \a      f       �T�f      j       \j      k       �T�                      @      y       U�      �       U	             U                      E      }       X�      �       X	              X                      N      }       Y�      �       Y	              Y                               W      \       0�_      }       P}      �       S�      �       P�      	       S	             P      [       Sf      g       S                       N      W       G�W      }       T�      �       T	              T                 +       2        0�                             +       2        0�2       @        S@       M        PM       U        S[       g        Sg       �        ]�       �        S                             +        1�+       X        \[       �        \                      �       	       U	             �U�             U                      �              T             �T�             T                      �              Q             �Q�             Q                      �              R             �R�             R                 �       �        0�                      �       �        X�       �        x��              p�                                     U        �       �U�                                  T                                    �        Q�       �        S�       �        �Q��       a       Sa      �       Q�      �       �Q�                                      )        0�)       8        P8       ;        p�;       ?        PB       �        Pa      }       P}      �       p��      �       P                             ?       	 x 0$0&�B       �       	 x 0$0&�a      �      	 x 0$0&�                   h       �        V�       a       V                    �       �        P$      0       P                        #       P                  M       �       V                 u       �        v�                     �       �        \�       a       \                    �       �        ]�       a       ]                    �       �        ^�       a       ^                    �       �        S�       �        s�                  G       �        S                          �      �       U�      �       �U��      �       U�      }       S}      ~       �U�                         �      �       u��      �       �U#��      �       u��      }       s�}      ~       �U#�                      #      &       q 7�&      K       QK      �       P                      �      �       U�      �       S�      �       �U�                  ;      ^       P                  E      n       T                          A      z       Uz      �       S�      �       �U��      �       S�      �       �U�                         A      z       u�z      �       s��      �       �U#��      �       s��      �       �U#�                                      U       ?        V?       B        �U�                                        T               T       >        S>       B        �TC%�                                      Q       A        \A       B        �Q�                      B       N        UN       ?       S?      A       �U�                  �       =       S                  �       $       P                           �      �       U�      �       �U��      �       U�      �       �U��      �       U�             �U�                    �             S             S                        �      �       P�      �       V�      	       v 1'�             v 1'�                      �      �       U�      �       S�      �       �U�                 �      �       V                      �      z       Sz      ~       U~             sH�      �       S                 �      �       S                      �      �       U�      �       �U��      �       U                  �      �       P                    �      �       P�      �       P                 �      �      ! p  $ &4$�ae     "� $ &2$u "                 �      �      ! p  $ &4$�ae     "� $ &2$u "                  �      �       V                  �      �       \                      	             P      c       Sc      n       s C%�                              N       p z �R      ]       p z �]      i       Qi      q       q C%�                          %       r s "�%      �       Y                          0      7       T7      9       t u �9      >       T>      E       XG      R       RR      T       r u �T      x       R                   �      �      
 �if     ��      �       P                  x      �       R                          �       P�      �       Q                              y      �       U�      x       Vx      }       �U�}      �       V�      �       �U��      �       V�      �       �U�                          |       U}      �       U                              v       Tv      |       t�}      �       T�      �       t�                      �      �       P�      �       S�             s C%�                        �      �       P�      �       p u ��      �       p u ��             Q             q C%�                       �      �       s p ��      |       X}      �       X�      �       X                        �      �       R�      �       r t ��      �       R�      �       R�      �       r t ��      1       R                    �              U      L       �U�                            �              T      C       VC      G       TG      H       �T�H      K       VK      L       �T�                     �              
 �if     �       B       SH      J       S                                 :        U:       �        V�       �        U�       �        V�       �        �U�                             *        T*       �        \�       �        �T�                         F       T        PT       a        Qa       e        q�e       p        Q�       �        v��       �        V                                     
 �if     �       �        S�       �        sx��       �        s��       �        sx�                                 P      �       S                    �      �       P�      �       S                      �      �       P�      F       SF      S       U                                                           0�      *       PK      U       PU      W       0�_      m       Um      �       V�      �       v��      �       U�      �       V�      �       0��      �       P             P      )       V)      ,       v�.      �       V�      �       0��      �       V�      �       v��      G       V                     <      S       \�      <       ]<      ?       }�                        m      �       UV      Z       PZ      n       U      5       U                  <      q       ]                  �      �       P                        A       _                      �
      �
       U�
      �
       V�
      �
       �U�                      �
      �
       P�
      �
       S�
      �
       P                      
      )
       U)
      ]
       V]
      ^
       �U�                  ,
      .
       P                  �	      �	       P                          m	      �	       S�	      �	       s��	      �	       v��	      �	       S�	      �	       V                  �	      �	       P                       �      �       Q�      �       q��      �       q2$p "�#��      �       Q                   a      m       ^m      �       ~j�                    �      �       ]�      j       ]                 �              ^                     �      �       Q�             ��      "       Q                                                  �      �       V�      �       v��      7       VK      W       V�      �       0��      �       _�      �       ��      �       _�      �       ^�      �       ~��      �       ^�      �       S�      �       s��      �       S�      �       U�      �       s��      �       S�      �       Q�      �       q��      �       q2$p "�#��      �       Q                                �      �       P�      �       p��      �       s 2$q "�#��      �       s 2$`�f     "�#��      �       R�             ��
      0       RV      [       1�[      h       P                      �      �       P�             \      .       V.      n       \                      7      =       P=      K       VW      �       V                    �      �       P�      �       \                   �      �       P�      �       s|�                  �      �       p��      �       S                  �      �       P�      u       ��                 @      �       0�                 �      �       \                    6      a       ^a      �       R                                  P             ��.      u       ��                  I      K       P                    �      �       P�      u       ��                    9      K       SW      [       S                                      P      �       ���      &       ��&      *       P*      u       ��                      M      Q       PQ      d       _k      {       _                      [      _       p�_      d       ~�k      n       ~�                     [      _       p  #>@s?@"�_      d       ~  #>@s?@"�k      n       ~  #>@s?@"�                  8      f       Q                   �      P       Vf      l       V                    "      *       p �f     ��*      8       Q                          �      )       U)      3       V3      E       UE      W       VW      X       �U�                    �      �       T�      �       v 2$`�f     "�t �                            -       P3      :       P:      E       v 3$@�f     "t "�0$0&�                           '       v 3$�f     "t "�
���'      -      5 �Tv 2$`�f     "� $ &1$v 3$�f     ""�
���3      E       v 3$�f     "t "�
���                        b      �       U�      �       P�      �       ^�      �       �U�                  �      �       S                       �      �       s��      [      
  3$s "#�[      ^      
  3$s "#$�^      `      
 3$s "#$�`      c      
  3$s "#�                  �      -       P                                    &       T&      V       RV      Y       r�[      `       Rc      �       _�      �       ��      �       _                        `       X                            #       R#      -       p �0$0&x "�-      `       U                     �      [       _[      ^       �`      c       _                  �      �       \                  �      �       ]                      N       �        U�       �        S�       b       �U�                      �       �        P�       U       VU      a       U                  o       [       ^                         �       �        ~��       5      
 s 3$~ "#�5      8      
 s 3$~ "#$�8      =      
 s3$~ "#$�=      O      
 s 3$~ "#�                  �       �        P                       �       �        y  $0 $+( ��       0       [0      3       {�5      =       [                  �       �        Y                    �       �        Q�       =       _                       �       �        0��       5       S5      8       s�=      O       S                  �       W       \                  �       Y       ]                          	        U	       N        X                          	        T	       N        Z                          	        R	       N        Y                               !        R!       #        x���#       +        R-       A        R                         ?        U                        K        x�                        ^
      o
       Uo
      �
       V�
      �
       �U��
      �
       U                      i
      o
       Uo
      �
       V�
      �
       �U�                  �
      �
       S                   p
      x
       p �f     ��x
      �
       Q                    �
      �
       P�
      �
       X                    �
      �
       P�
      ;       Y                     �
      �
       X�f     �x "
@y ��
      �
       U      ;       X                       ;       Z                    k
      �
       U�
      �
       �U�                      k
      �
       T�
      �
       R�
      �
       �T�                  j      �       P                        q      {       [�      �       Q�      �       U�      �       q@��      �       Q                            �      �       0��      �       S�      �       sx��      	       S	      1	       S1	      6	       sx�6	      D	       S                           q      {       0�L	      k	       Sk	      p	       sx�p	      ~	       S�	      �	       S�	      �	       sx��	      a
       S                        �      �       P�      	       V	      	       P	      L	       VL	      L	       PL	      �	       V�	      �	       P�	      b
       V                  e      i       U                           �      �       Q�      �       q��      �       Q�      �       Q�      �       q��      �       Q                   �      V       P�      �       P                        �       R                   ;      R       p J%�R      f       X                   ;      V      	 p 4%
��\      _       Q                     ;      K       TK      _       t~�s      �       T                           T       UT      �       u��      �       U                 ;      V       p 4%
�p J%!�                   %      d       P�      �       P                  6      �       Q                  I      �       U                    Q      [       T[      �       t��      �       T                 Q      d       p 4%
�p J%!�                   Q      b       p J%�b      t       X                   Q      d      	 p 4%
��j      m       R                     A      F       0�F      �       p�~��      �       p�~�                      =      A       q t �A      �       V�             v�      $       V                      �      �       X�             x q "�            	 x q "#��      $       x q "�                      �      �       U�             u q "�            	 u q "#��      $       u q "�                    �      �       P�      �       R      $       P                 �      $       T                    Y      �       S�      $       s�                            �       q t ��      �       S�      '       s�'      ,       S                    �             Q      '       q�}�'      ,       Q                     �      �       P�      �       R'      ,       P                 �      ,       T                      �      �       q t ��      W       VW      j       v�j      o       V                    �      ^       R^      j       r�}�j      o       R                           d       Pd      j       p�}�j      o       P                              	 p�f                        �      �       S�              s�                      �      �       q t ��      G       SG      S       s�S      X       S                          M       PM      S       p�}�S      X       P                            	 p�f                           �       �        q t ��       R       SR      s       s�s             S                      B      G       TG      s       t q "�s      z      	 t q "#��z             t q "�                      E      G       RG      s       r q "�s      z      	 r q "#��z             r q "�                    E      U       PU      X       Us             P                 E             X                            &       Q&      ?       q�?      G       ��f     �1$�                                     q t �       �        S�       �        s��       �        S                    u       �        Q�       �        q�}��       �        Q                     {       �        P�       �        R�       �        P                 u       �        T                    	      	       U	      J	       �U�                   �      �       Q�      �       q�                      �             U      4       V4      D       �U�                      �             T      8       \8      D       �T�                        /       S                  &      -       P                          %       P-      2       P                  �      �       T�      �       t �                                 C      E       0�E      Q       PQ      T       p�V      ]       P]      �       S�      �       s��      �       S�      �       s��      �       S                                  0�      B       TB      E       t�                           -       t 
@r 	�x "�-      2       p  $0 $+( �2      c      $ q { q  $O $,(  $0 $+( �                         V       XV      c       x�                 C      X       0�                     X      ]       0�]      �       v��      �       V                     l      r       p <&	�} "��      �       p  $0 $+( ��      �      # r Or  $O $,(  $0 $+( �                   X      �       ]�      �       }�                    l      l       Pl      r       p <&�r      u       P                  �      �       Q                        �      �       P�      �       p��      �       u��      �       P                            u      w       P~      �       P�      �       P�      �       Q�      �       P�      �       | <�f     "                  Q      Q       PQ      9       S                    �      �       U�      3       �U�                        $       P                	   �      �       u �f     �@J$"��      �       �U�f     �@J$"�                  �      1       S                    �      �       P�      2       V                  �             P                        E      |       U|      �       �U��      �       U�      �       �U�                    E      S       TS      �       �T�                      a      x       Px      �       S�      �       P                          j      v       Sv      x       Qx      �       P�      �       S�      �      	 t r 'r �                    �      �       P�      �       P                      0      8       U8      D      	 zg     D      E       �U�                      0      @       T@      D      	 zg     D      E       �T�                    0      D       QD      E       �Q�                    0      D       RD      E       �R�                                          %      ;       U;      _       U_      c       Tr      y       U�      �       U�      �       T�      �       U�      �       U�      �       R�      �       R�             R             R/      0       U                                        %      >       T>      c       Xr      y       X�      �       X�      �       Q�      �       Q�      �       X�      �       X�      �       X�             Q             Q/      0       X                      �       �        U�       $       �U�$      %       U                      �       �        T�       $       �T�$      %       T                    �       �        Q�       %       �Q�                    �       �        R$      %       R                   �       	       X$      %       X                                �       �        p r ��       �        P�       �        �Q#�r ��       �        P�       �        S�       �        P�              S$      %       �Q#�r �                    �       	       Q$      %       Q                    �       �        P�       	       P                      �       �        T�       �        T�              V                                 P             \                               P                             w        Uw       �        �U��       �        U                             ^        T^       �        �T��       �        T                               �        Q�       �        S�       �        �Q��       �        Q                  [       �        R                    g       |        T|       �        V                    �       �        P�       �        \                  �       �        P                  �      �       S                    �      �       P�      �       p  $? $-( �                        �      (       V(      +       v��      �       ]�      �       U�      �       ]                 �      �       ^                               T                  J      �       V                      @      d       Ud      �       ^�      �       ���#�                           @      d       Tg      �       ]�      �       U�      �       _�      �       ]�      �       _                            @      d       Qd      �       S�      �       S�      �       U�      �       S�      �       T                        @      d       Rd      �       \�      �       Q�      �       q��      �       Q                        @      d       Xd      �       V�      �       X�      �       x��      �       X                          �              U       '       �U�'      1       X1      <       U<      @       X                        �             Q      1       x1      <       Q<      @       �Q�                 �      �       P                 �      �       R                  �      @       Y                 �      �       X                   �      �       P1      <       P                    '      J       UJ      �       ]                      '      �       T�      �       \�      �       �T�                    '      J       QJ      �       V                     J      Q      
  �g     �Q      �       S�      �       P                       �      �       0��      �       P�      �       p��      �       P                  �             S                             <        U<       �       ]�      �       �U�                             7        T7       �       V�      �       �T�                             5        Q5       �       \�      �       �Q�                  �       �       ^                          }       �        P�       �        S�       �        S�       �        U�       J       S                      �       �        P�              Q      �       ��                  J      J       SJ      V       s ��������-( �                        -      g       Ug      �       S�      �       �U��      �       U                              -      b       Tb      E       \E      P       PP      t       �T�t      x       \x      �       �T��      �       T                    �      �       P�      �       ��                      �      �       Q�      �       V�      �       Q                         �      �       p (�i     ���      �      " p (�i     � $@J$ $-( ��      �      +  �i     �(�i     � $@J$ $-( ��	      �	       P�	      �	       q p ��	      �	       P�	      �	       p ����@J$����-( �                  i
      �
       P                                 P      &       p ����/����-( �&      P       r <&����/����-( �                    P      7       S7      ?       s�                  �      $       \                    �      ,       ^m      �       S                        $       ]                    o      �       X�      �       T                   o      �       T�      �       Q                                �        U�              �U�             U             �U�                            D       TD             �T�                                      Q              V             �Q�                    �      �       P�      �       p ����/����-( ��      �       t <&����/����-( �                    �      �       p}��      �       U                  V       �        P                  ?              S                  q      �       S                      h      j       S�      �       S�      �       S                        ?      x       Ux      C       \C      I       UI      J       �U�                  x      A       V                	                          ?      A       uP      h       Ph      k       p�m      t       PD      h       Th      k       t�u      �       T�      �       t��      �       T�      �       t��      �       |�              P       #       p�%      ?       P                  �      �       S                  �      �       ]                    �      �       Q�             Q                    �      �       P�             P                                /       P/      2       p 	��2      4       P<      A       Pm      u       P�      �       P                   �             R      <       r�<      ?       R                    �      �       R�      ?       Y                        �      �       P�      �       p���      �       P�      �       P�             Q                  �      >       P                     �      �       �����      �       U�             U                   .      <       0�<      U       1�                  �
             P                           .      7       s��7      ;       U;      <       s��<      M       s��M      R       US      T       s��                      �      �       U�      �
       ]�
      �
       �U�                 a	      �	       S                  �	      �
       _                    �	      �	       q��	      �	       Q                  	      a	       S                    K	      X	       PX	      a	       } #�
�����Ls"�                  [	      �
      	 ~ 0$0&�                 [	      �
       | ��                 �	      �
       W                      o      �       U�      �       �U��      �       U                  �      �       S                  �      �       P                      �      �       U�      n       _n      o       �U�                  �      L       S                  �      �       ]                                     P             \L      P       p �P      S       s �                          1       p �Q      Z       P                 S      0       S                          -       \-      1       T                    <      @       P@      H       V                  #      `       \                    O      Q       t�Q      �       T                  �      	       ]                  �             \                    �      �       ^�      `       ^                  �      �       P                    �             P      `       ��                  H      H       VH      N       v  $/ $-( �                    l      s       Ps      `       S                  �      �       P                      �      �       P�      �       p ��      �       P                      �      �       U�      �       S�      �       �U�                    �      �       T�      �       �T�                    �      �       Q�      �       �Q�                   �      �       }  $ &2$v "#� $ &v "��      �       | @& $ &2$v "#� $ &v "�                       }      �       | @&��      �       ]�      �       | @&��      �       ]                 Z      �       \                    �      �       P�      �       V                  �      �       U�      �       S                            %       Q%      /       r��|�/      y       p ��i     ��i     �"�                             %       t q "�%      ,      
 r t "
���,      /       s����i     �r��|"�/      8      / s����i     �p ��i     ��i     �""�                  �      �       V                    �      �       U�      �       �U�                     �      �       0��      �       P�      �       p�                        B      {       U{      �       V�      �       �U��      �       U                
   B      E       UE      T       P                       �      �       0��      �       S�      �       s��      �       S                 �      �       \                        &      A       TA      J       ��f      m       t 8$8&A�m      |       t� 8$8&A��      I       ]                           )      A       QA      J       ��f      x       p�8$8&0�x      |       Q�             y�      .       Y                    �      �       ~��      �       �                    �      �       p��      �       ���#�                  J      R       P                                  )        U)       �        \�       �        �U��              \      B       �U�                              $        T$       9       V9      B       �T�                            /        Q/       �        ^�       6       ~�                              /        R/       =       ]=      B       �R�                   �       �        P�       �        p�                      P      Z       UZ      k       Xk      l       �U�                  P      ^       T                    2      J       UJ      P       �U�                    2      8       T8      P       �T�                      9      K       UK      /       \/      2       �U�                        9      G       TG      ,       S,      -       vh�-      2       �T�                        U      ^       P^      a       Va      a       sf      q       Pq      �      
 s�6$q "�                  a      �       V                       U      ^       p 6$�^      c       Pc      n       s�6$�n      �       ]                               �      �       V�      �       s��      �       s��      �       s��      �       s��      �       s��      �       s��      �       s��             s �             s!�             s"�             s#�             s$�             s%�             s&�             s'�             s(�             s)�             s*�             s+�      ,       s,�,      -       v�-      2       �T#,�                      W      x       Ux      1       S1      9       �U�                             W      t       Tt      �       V�      �       T�      �       V�      �      	 v | "} �             v q "�      *       v q "#�*      0       v q "�                                W      x       Qx      �       \�      �       Q�      �       \�      �       ]�      �       }� ��             ]      *       | q �*      .       | q #�                            �        U�       +       ��~                            >        T>       D        t�D       K        t}�K       Q        t~�Q       W        t�W       �        T                                                                                             P        �        u �       �        ��~�       $       R$      S       ��~�2# $��������%!�S      {       X�      �       X�      '       T@      t       T�      �       U�      �       U�      �       S�      s       S{      �       S�      �       S�      B       Sd      �       S	      >       Sa             S      a       Qa      g       X|      �       Q3	      �	       X�	      �	       P�	      i
       X�
      �
       P�
      �       P�             U      !       Q;      �       U�      O       YY             Y      j       ]v      \       ]c      �       ]�      T       ]d      �       ]�      �       T                                                                            $       '        P'       �        u�       �        ��~#�       �        U�              X      1       ���2# $��������%!�1      \       T\      p      ���~�2# $��������%!��~���~�'�����~�'��~�5$��������# %!"���"z "#���2# $��������%!'���2# $��������%!��~�'��~���~�'��~���~�'�����~�'��~�5$��������# %!"���"z "#���5$��������# %!"��~�"{ "#�����~�2# $��������%!'���2# $��������%!��~�2# $��������%!'��~���~�'�����~�'��~�5$��������# %!"���"z "#������2# $��������%!'���2# $��������%!��~�'��~���~�'��~���~�'�����~�'��~�5$��������# %!"���"z "#���5$��������# %!"��~�"{ "#���5$��������# %!"��~�"s "#���5$��������# %!"���2# $��������%!"v "#����p      �       T�      �      ���~�2# $��������%!��~���~�'�����~�'��~�5$��������# %!"���"z "#���2# $��������%!'���2# $��������%!��~�'��~���~�'��~���~�'�����~�'��~�5$��������# %!"���"z "#���5$��������# %!"��~�"{ "#�����~�2# $��������%!'���2# $��������%!��~�2# $��������%!'��~���~�'�����~�'��~�5$��������# %!"���"z "#������2# $��������%!'���2# $��������%!��~�'��~���~�'��~���~�'�����~�'��~�5$��������# %!"���"z "#���5$��������# %!"��~�"{ "#���5$��������# %!"��~�"s "#���5$��������# %!"���2# $��������%!"v "#���2# $��������%!��             U      U       U�      �       P�      Q       Pe      �       P�      B       PP      �       V�      p       Vx      �       V      �       V�             Y+      �       Y�             R             P2      �       R		      ^	       R^	      `	       Q	      K
       YK
      �
       Q�
      p       Qx      �       X�      �       X�             ["      7       [R      2       [?      �       [�              [+      �       [�      �       R                                                                          +       .        P.       �        u�              ��~#      P       UP      S      b���2# $��������%!��~�2# $��������%!'��~���~�'�����~�'��~�5$��������# %!"���"z "#������2# $��������%!'���2# $��������%!��~�'��~���~�'��~���~�'�����~�'��~�5$��������# %!"���"z "#���5$��������# %!"��~�"{ "#���5$��������# %!"��~�"s "#����S      �       U�      �      z���2# $��������%!��~�2# $��������%!'��~���~�'�����~�'��~�5$��������# %!"���"z "#������2# $��������%!'���2# $��������%!��~�'��~���~�'��~���~�'�����~�'��~�5$��������# %!"���"z "#���5$��������# %!"��~�"{ "#���5$��������# %!"��~�"s "#���2# $��������%!��      �       P�      1       Pc      �       Q�             Q'      �       Q�             Q      ]       \{      /       \7      �       \�      j       \�      �       Z	      n       Z�      �       T      �       T�      	       T	      	       X3	      �	       T�	      l
       Rl
      n
       P�
      0       R8      �       Y�      +       Ya      �       V�      �       V�      �       U      �       U�             Z      �       Z�      �       S�      �       S                                                                                2       5        P5       �        u�       �        ��~#�              P      1      � ���2# $��������%!��~�'��~���~�'��~���~�'�����~�'��~�5$��������# %!"���"z "#���5$��������# %!"��~�"{ "#����1      f       Pf      �      � ���2# $��������%!��~�'��~���~�'��~���~�'�����~�'��~�5$��������# %!"���"z "#���5$��������# %!"��~�"{ "#���2# $��������%!��      �       Q�             Q@      �       R�      T       Re      �       R�      F       ]P      �       ]�      e       ]x      W       ]d      �       ]�      Y       ]a      �       U�      ^       U|      �       U�      �       X		      �	       U�	      
       P
       
       QM
      O
       PO
      �
       T�
      [       Z[      `       Rx      ;       Z;      �       R�      Q       RY      �       X�      o       Xv      �       V�      T       Vc      �       V�      P       Vd      �       U                                                                                9       >        P>       �        u�       �        ��~#�       �        Q�             E ��~���~�'�����~�'��~�5$��������# %!"���"z "#����      E       QE      p      ] ��~���~�'�����~�'��~�5$��������# %!"���"z "#���2# $��������%!�p      �       R�      �       R      K       Xc      �       X�             T'      �       T�             [      �       [�      $       [7             [      T       [�             [+      �       X�             X2      �       P�      V	       P	      �	       Q�	      �	       U�	      �
       U�
             [              T8      �       [�      J       TJ      L       Qa             T"      s       T�      J       TR      �       \�      7       \?      �       \�             \+      �       X�      �       Q                                                                                                                                                                                                           e      ~       v } '���'z '�~      �       X�      �       v } '���'z '��      �       | ~ '���'y '��      �       U�      �       | ~ '���'y '��      �       } ���'���'��~�'��      �       T�      �       } ���'���'��~�'��      �       ������'���'��~�'��             ~  '�@�'x '�             R             ~  '�@�'x '�      4       ������'�D�'u '�4      9       Q9      P       ������'�D�'u '�P      c        w �'z 't '�c      l       ���w �'z 't '�l      q       Pq      {       ���w �'z 't '�{      �       ������'y 'r '��      �       ^�      �       ������'y 'r '��      �       w ����'��~�'q '��      �       ^�      �       w ����'��~�'q '��             ������'x 'p '�             ^      7       ������'x 'p '�7      I       ����@�'u '��~�'�I      O       ^O      x       ����@�'u '��~�'�x      �       ����D�'t '��~�'��      �       ^�      �       ����D�'t '��~�'��      �       �@�z 'r '��~�'��      �      > ������'���'���'1$��������# %!�@�'r '��~�'��      �       ^�            > ������'���'���'1$��������# %!�@�'r '��~�'�      !       �D�y 'q '��~�'�!      .      = ������'���'�@�'1$��������# %!�D�'q '��~�'�.      1       ^1      d      = ������'���'�@�'1$��������# %!�D�'q '��~�'��      �       ��~�u '��~�'��~�'��      �       V�      �       ��~�u '��~�'��~�'��      �      k ������'���'�@�'1$��������# %!���'���'���'1$��������# %!��~�'��~�'��~�'��      	      � ������'w �'�D�'1$��������# %!������'���'�@�'1$��������# %!���'���'���'1$��������# %!'��~�'��~�'�2      A       ��~���~�'��~�' '�A      I      � ������'���'�@�'1$��������# %!������'���'���'1$��������# %!���'���'���'1$��������# %!���'���'�@�'1$��������# %!'���'���'1$��������# %!��~�'��~�' '�I      O       XO      U       _U      |      � ������'���'�@�'1$��������# %!������'���'���'1$��������# %!���'���'���'1$��������# %!���'���'�@�'1$��������# %!'���'���'1$��������# %!��~�'��~�'��~�'�|      �       ��~���~�'��~�'{ '��      �       ^�      	       ��~���~�'| 's '�	      		      5������'���'���'1$��������# %!���'���'���'1$��������# %!������'���'���'1$��������# %!������'w �'�D�'1$��������# %!���'���'���'1$��������# %!'���'w �'1$��������# %!'���'���'1$��������# %!��~�'| 's '�		      3	       ��~���~�'v ' '�3	      B	       ��~���~�'} '��~�'�B	      D	       QD	      	       ��~���~�'} '��~�'�	      �	       ��~���~�'��~�'��~�'��	      �	       R�	      �	       ��~���~�'��~�'��~�'��	      
       ��~���~�'s '{ '�
      #
       Z#
      M
       ��~���~�'s '{ '�M
      \
       ��~�| ' '��~�'�\
      a
       Za
      �
       ��~�| ' '��~�'��
      �
       ��~�v '��~�'��~�'��
      �
       | } '��~�'��~�'��
      �
       X�
      �
       | } '��~�'��~�'��
             v ��~�'��~�'��~�'�             U      8       v ��~�'��~�'��~�'�8      I       } ��~�'��~�'~ '�I      N       TN      x       } ��~�'��~�'~ '�x      �       ��~�s '��~�'��~�'��      �       R�      �       ��~�s '��~�'��~�'��      �      Q������'���'���'1$��������# %!���'���'���'1$��������# %!���'���'�@�'1$��������# %!������'���'���'1$��������# %!������'w �'�D�'1$��������# %!���'���'���'1$��������# %!'���'w �'1$��������# %!'������'���'���'1$��������# %!������'���'���'1$��������# %!���'���'���'1$��������# %!���'���'�@�'1$��������# %!'������'���'���'1$��������# %!���'���'���'1$��������# %!������'���'���'1$��������# %!������'w �'�D�'1$��������# %!���'���'���'1$��������# %!'���'w �'1$��������# %!'���'���'1$��������# %!'�@�'1$��������# %!'| '1$��������# %!s '��~�'��~�'��      �       ��~� '��~�'��~�'��      �       P�      �       ��~� '��~�'��~�'�a      u       ��~���~�'~ 'p '�u      z       Yz             ��~���~�'~ 'p '��      �       ��~���~�'��~�'s '��      �       X�      �       ��~���~�'��~�'s '��              ��~���~�'��~�' '�       	       U	             ��~���~�'��~�' '�"      2       ��~���~�'��~�'��~�'�2      6       Q6      :       ��~���~�'��~�'��~�'�Y      n       ��~���~�'��~�'z '�n      u       Ru      y       ��~���~�'��~�'z '��      �       ��~�~ 's '��~�'��      �       R�      �       ��~�~ 's '��~�'�             ��~���~�' '��~�'�              Z       F       ��~���~�' '��~�'�R      v       ��~�~ '��~�'��~�'�v      �       ��~���~�'��~�'��~�'��      �       X�      �       ��~���~�'��~�'��~�'��      �       ��~���~�'��~�'��~�'��      �       U�      �       ��~���~�'��~�'��~�'�      +       ��~�s '��~�'x '�+      4       R4      ?       ��~�s '��~�'x '��      �       ��~���~�'y 'p '��      �       Y�             ��~���~�'x 'q '�      
      ? ��~���~�'��~�'��~�'1$��������# %!��~�'��~�'q '�
             Q+      8       ��~���~�'u 'z '�8      >      ? ��~���~�'��~�'��~�'1$��������# %!��~�'��~�'z '�>      J       Zd      �       ��~���~�'t 'y '��      �       T�      �       ��~���~�'r 'q '��      �       R�      �       ��~���~�'p 'z '��             Z                 9       >        0�                       9       >        ���>       H        PH       ]        p|�]       k        P                              	        U	       C        SC       D        �U�                        �      ,       U,      �       S�      �       �U��      �       U                      �      7       T7      �       �T��      �       T                        �       |  0$0&�                  $      �       V                 $      �      	 } 0$0&�                 $      �      	 ~ 0$0&�                        �      /       U/      �       S�      �       �U��      �       U                      �      k       Tk      �       �T��      �       T                 S      �       ]                   S      k       Xk      q       �L                  M      �       \                  S      �       V                        �      �       U�      �       S�      �       U�      �       �U�                        �      �       T�      �       V�      �       T�      �       �T�                 �      �       3�                 �      �       Y                 �      �       X                 �      �       R                 �      �       Q                 �      �       T                 �      �       U                      z      �       U�      �       �U��      �       U                      z      �       T�      �       �T��      �       T                          9       �        U�       ^       V^      k       �U�k      q       Vq      z       �U�                    9       �        T�       z       �T�                         X       �        ^�              S             0�      +       S;      E       S                    f       f       _k      y       _                    k       �        X�       �        ��                     k       b       ]b      j       u�k      u       ]                   o       d       ~  $0-��k      w       ~  $0-��                   X      \       0�\      �       S                
     x      z       0��      �       0��      �       1��      �       2��      �       3�                    s      {       U{      �       �U�                      s      {       T{      �       S�      �       �T�                                    U               �U�                              	        T	               S               �T�                             $        U$       k       Sk      s       �U�                                   $        0�$       i        Vi       m        R�       �        V�       	       VS      0       V0      4       R4      E       v�E      l       V                       S      Y       0�Y      r       ]r      v       Xv      �       }��      p       ]                           S      S       0�S      Y       v 3$�Y      r       v 3$} "�r      v       v 3$x "�v      �      
 v 3$} "1��      �       v 3$#��      �       v 3$#��             v 3$#�      0       v 3$#�0      4       r 3$#�4      E       v3$#�Z      f       )�f      s       *�                    �      �       U�      �       �U�                  �      �       T                        �      �       U�      �       S�      �       T�      �       �U�                       V      b       0�b      n       1�n      z       2�z      �       3�                                       S+      6       SQ      |       S|      �      	 4f     �      �       S                      �             S             sy�             S                       �      �       <q 6&��      �       <r 6&��      �      	 <p<�6&��      �       Q                                         0�      (       P(      +       p�+      5       q~��      �       0��      �       Q�      �       q�                  B	      f	       X                    	      	       P(	      4	       P                    "	      (	       P*	      f	       U                    6      E       RE      P       1�P      v       R                  �      �       R                        �      I       UI      �       S�      �       �U��      �       U                              	      	       0�	      	       1�	      	       2�	      0       3�0      5       4�r      r       0�r      r       1�r      r       2�r      �       3��      �       0��      �       1��      �       2��      �       3��      �       4��      �       5��      �       6��      !       V!      $       v�                                   p q "@�!      )       �^�8$8&p "0�@      D       �^�8$8&p "0�                         +       1�.      E       T                    $      +       Q1      �       Q                          �      �       U�      �       U�      �       T�      �       U�      �       p�                          �      �       T�      �       V�      �       T�      ^       V^      _       �T�                   �      �       0��      ]       S                  C      P       P                    �      �       U�      �       �U�                      �      �       U�      �       S�      �      	 t%f                             h      y       Uy      �       S�      �       U�      �       �U�                      �      �       U�      c       \c      h       �U�                  3      I       P                          �      S       SS      V       s�V      [       }�[      `       S`      e       ]                  �      [       ^                  �      [       V                      �      �       U�      P       \P      S       �U�                      �      �       T�      �       S�      S       �T�                      �      �       U�      P       \P      S       �U�                        O       P                       H       ]                b             \                          b      o       0�o      �       ]�      �       P�      �       ]�      �       P�             ]                               P                      D       R        UR       W       ]W      X       �U�                    D       _        T_       X       �T�                      D       �        Q�       P       SP      X       �Q�                      D       �        R�       P       \P      X       �R�                    �       	       V	             v  $�C$ $-( �1      F       V                    o       �        P�       �        u { u { O&'u { O&�                  �       �        X                  �       �        P�       �        p C%�                      X      y       Uy      ~       �U�~      �       U                     X      g       0�g      }       P~      �       P                       _      f       0�f      �       S�      �       s��      �       S                    �      �       U�      �       U                           $        U$       D        �U�                 5       B        0�                         C        S                      �      �       U�      8       V8      =       �U�                      �      �       T�      2       S2      =       �T�                   �      �       Q�      	       Q	             1�                                    U       )        �U�                                    T       )        �T�                          (        P                          �	      �	       U�	      �
       S�
      d       �U�d      i       Si      s       �U�                    �	      �	       P�	      s       ��                      �	      
       P
      _       _d      r       _                        
      
       P
      Y       \Y      d       Rd      l       \                      !
      %
       P%
      ]       ^d      p       ^                          =
      �
       P�
             V      ,       R,      R       Vd      s       P                      8
      <
       P<
      [       ]d      n       ]                 �
      d       ��                 �
      d       ?�                   �
      �
       s r ��
      �
       S                 �
      d       (�                    �
      �
       P�
      d       X                      A	      L	       UL	      �	       V�	      �	       �U�                   A	      L	       0�L	      �	       S                      4      `       U`      4	       V4	      A	       �U�                          4      L       TL      �       ]�      �       } p "��      �       } p "#��      �       } p "��      �       } p "#��      	       } p "�                      4      S       QS      6	       \6	      A	       �Q�                      4      m       Rm      <	       _<	      A	       �R�                        4      m       Xm      	       ��	      	       X	      	       x p "�	      	       x p "#�	      *	       x p "�                           �      �       0��      �       P�      �       p��      	       P	      	       0�	      	       P	      	       p�                 	      	      	 q s #��                      {      �       P�      3	       S3	      @	       U                           �      �       Q�      �       q��      �       Q�      �       q��      �       q��      �       Q�      	       q�	      	       q p "#�	      	       q p "#�	      	       q p "#�	      &	      
 q p "
 �                      
             U             T             �U�                    �      �       U�      
       Z                    �      �       T�      
       Y                      �      �       Q�             S      
       �Q�                    �      �       R�      
       [                  �      �       U�      �       �U�                    �      �       T�      �       �T�                     �      �       T�      �      
 p 
@t "��      �      
 p
@t "��      �      
 p 
@t "�                   �      �       P�      �       P                          �       T�      �       �T�                    �      �       T�      �       t p "��      �       t p "#��      �       t p "�                     �      �       P�      �       p��      �       P                    E      [       U[             �U�                    E      K       TK             �T�                  ^             U                        f      j       u p "�j      q       p u "#�q      s       p u "�s      z       u p "�z      ~      
 u p "
@�                      f      n       Pn      q       p�s      ~       P                   ^      `       0�`             T                      �      �       U�      D       ^D      E       �U�                        �      �       T�             S             T      E       �T�                      �      �       Q�      >       V>      E       �Q�                    �      �       R�      B       ]                        �      �       X�      :       \:      <       T<      @       \                            5       S5      7       U7      :       s�}�:      =       S                     �      �       U�      �       u p ��      �       U�             V                      �      �       T�      �       �T��      �       S                      �      �       Q�      �       \�      �       �Q�                   6      6       r���6      ^      
 v  ~ �"�l      w      
 v  ~ �"�                      �             0�      w       Qw      z       q�|      �       Q                        |       R                                       T      w       [w      z       t q "#�z      |       t q "�|      �       [                    3      6       ]6      c       } u "�c      j      	 } u "#��j      w       } u "�                         6       r�6      V       r v "#�V      ^       r v "#�^      u       r v "#�                                        Y      w       Sw      z       y q "#�z      |       y q "�|      ~       S~      �       y q "�                    6      6       P6      V       p u "�V      j      	 p u "#��j      p       p u "�                       �       Z                     �      �       U�      �       u p ��      �       U�             \                      �      �       T�      �       �T��             S                      �      �       Q�      �       V�      �       �Q�                 C      �       U                      �             0�      �       T�      �       t��      �       T                  *      �       Q                                      S      �       Y�      �       s t "#��      �       s t "��      �       Y                    C      W       PW      t       p�}�t      z       P                     1      @       q�@      J       ZJ      Z       z�Z      �       Z                       �       X                      �             U             �U�      H       \                        �             T             �T�      "       S8      H       S                          �             Q      8       V8      :       Q:      �       V�      �       �Q�                 v      �       Z                           8       0�H      K       t�O      �       T                    H      K       R\      �       R                      6      8       SH      K       s t "#�O      �       Y                    v      �       P�      �       p�}��      �       P                    s      �       U�      �       u��      �       U                   6      8       XH      �       X                     (      ;       U;      =       u p �=      e       Ue      �       \                      (      5       T5      ;       �T�;      r       S                      (      k       Qk      �       V�      �       �Q�                 �      �       U                      l      �       0��      �       T�      �       t��      �       T                  �      �       Q                         �      �       S�      �       Y�      �       s t "#��      �       s t "��      �       Y                    �      �       P�      �       p�}��      �       P                     �      �       q��      �       Z�      �       z��      �       Z                 �      �       X                    #      '       U'      (       �U�                    #      '       T'      (       �T�                    #      '       Q'      (       �Q�                     -      B       UB      L       �U�L      �       \                        -      :       T:      @       �T�@      �       S�      �       T                          -      Q       QQ      X       VX      Z       QZ              V       #       �Q�                   �      �       p����            
 r  z �"�
            
 r  z �"�                    �      �       0��             T             t�                  �             P                       �      �       S�             Y             s t "#�             s t "�                     �      �       Q�            
 r 
@q "�            
 r
@q "�
            
 r 
@q "�                   �      �       p��      �       p r "#��             p r "#�             p r "#�                 �             X                     +      @       U@      J       �U�J      �       \                        +      8       T8      >       �T�>      �       S�      �       T                          +      O       QO      _       V_      a       Qa      *       V*      -       �Q�                   �      �       p����            
 t  y �"�      #      
 t  y �"�                    �      �       0��      #       R#      &       r�                  �      (       P                       �      �       S�      #       X#      &       s r "#�&      (       s r "�                     �      �       Q�            
 t 
@q "�            
 t
@q "�            
 t 
@q "�                   �      �       p��             p t "#�             p t "#�      !       p t "#�                 �      (       U                      K       �        U�               ^       #       �U�                      K       �        T�              V      #       �T�                    K       �        Q�       #       ��                      K       �        R�              \      #       �R�                    K       �        X�              ]                      K       �        Y�       "       _"      #       �Y�                      �              Q             T             q�}�      #       Q                 �       #       Y                                )        U)       @        S@       J        �U�J       K        U                                  !        T!       .        Q.       A        VA       J        �T�J       K        T                                        Q       C        \C       J        �Q�J       K        Q                                .        R.       E        ]E       J        �R�J       K        R                      $       .        R.       E        ]E       J        �R�                    $       C        \C       J        �Q�                      $       )        U)       @        S@       J        �U�                    �      �       U�      �       �U�                    S      [       U[      e       �U�                      S      [       T[      d       Sd      e       �T�                                    U               �U�                              	        T	               S               �T�                             /        U/       I       SI      S       �U�                                     /       b        Vt       y        0�y       �        V             0�      R       YR      _       \_      k       Yk      n       |�t      |       Y|      �       V�      �       V�      �       r�                      �       t       Vt      w       v�w      |       �                                 Z      |       ^                     �      �       0��      �       T�      �       t�                  �             P                        �      �       P�      �       S�      y       vN�~      �       vN�                   �      o       So      r       s�                                  �      �       \�             |� �             U             |� �      %       |��%      *       U*      /       |��/      >       |��>      C       UC      H       |��H      `       |��`      j       Uj      o       |��                  �      �       ]                  i             V                         j      u       0�u      �       X�      �       x��      �       X�      �       x�                  �      �       P                              c       U�      �       U      _       U�      �       Z                   �             X             x�                     @      �       S�      �       s�             0�"      ~       S~      �       s�                     0      0       R�@      �       ^�      �       s (#z�"      5       R�5      Y       v :#R�Y      ]       v :#z�                     0      0       D�@      �       ]�      �       s !#e�	             N�"      ~       \~      �       s !#o�                          �       ]�      �       ~��                         �
      �
       0�      E       UE      U       u��      A       UA      Z       u�                  �      ^       Y                     &
      8
       0�8
      J
       QJ
      M
       q�                   &
      8
       0�8
      S
       PS
      W
       p u  $ &#2$r "#��                         �	      �	       0��	      �	       V�	      �	       U�	      �	       v��	      
       V                  �	      
       S                          ?      �       U�      �       Y�      �       ���      �       Y�             S                      ?      �       T�             _             �T�                                ?      t       Qt      �       \�      �       Q�      �       \�      �       Q�      �       P�      �       ���      �       Q                          ?      t       Rt      w       Vw      y       v�y      �       V�      �       R�      �       S                  c             ]                 }      �       |  $0-��                  t      }       P                      �      �       U�      ^       R^      f       �U�                    �             T      f       �T�                 �             0�      _       1�                            �      �       Y�             u q�0$0&�             u t #�0$0&�             u �T#�0$0&�      9       X9      P       u q�0$0&�                     �             p q�0$0&�             p t #�0$0&�             p �T#�0$0&�      P       p q�0$0&�                                 �      �       q �0$0&y "��      �       X�      �       q �0$0&y "��             q �0$0&q�0$0&u "�             t �0$0&t #�0$0&u "�             �T�0$0&�T#�0$0&u "�      %       q �0$0&x "�%      6       T6      9       q �0$0&x "�9      P       q �0$0&q�0$0&u "�                     �             q�0$0&q�0$0&p "�             t #�0$0&t #�0$0&p "�            ! �T#�0$0&�T#�0$0&p "�             �T#�0$0&q�0$0&p "�      P       q�0$0&q�0$0&p "�                     5             2�      �       r�0$0&54#��      �       q�0$0&54#�                   x      �       2��      
      3 �'f     #� $ &3$0&f     "#�0$0&54#�
      )       2�                      �      �       V�             v�             V                  �             S                          -      �       \�      �       T�      �       \�      �       |��      �       T                  T      �       S                             7       S7      :       s�<      =       S                        6       P                                -       U-      9       S9      @       U@      A       �U�A      B       U                                -       T-      :       V:      @       T@      A       �T�A      B       T                                #       Q#      <       \<      @       Q@      A       �Q�A      B       Q                      )      <       \<      @       Q@      A       �Q�                        )      -       T-      :       V:      @       T@      A       �T�                        )      -       U-      9       S9      @       U@      A       �U�                                B      m       Um      �       V�      �       P�      �       V�      �       U�      �       �U��      �       V�      �       U                              B      m       Tm      �       ]�      �       T�      �       �T��      �       ]�      �       �T��      �       T                                B      m       Qm      �       \�      �       Q�      �       \�      �       �Q��      �       \�      �       �Q��      �       Q                     m      �       S�      �       S�      �       S                 m      �       | s <�                      �      �       Q�      �       \�      �       �Q�                    �      �       U�      �       �U�                  �      �       U                                    U              ��~                     ,       �        V�       �        v��       �        V                  O       �        S                                  O       \        ��~�\       e        Ue       �        ��~��       �        U�       �        ��~��       �        U�       �        ��~��       �        U�       �        ��~�                 j       �        ]                      |       �        P�       �        T�       �        P                    !       &        U&       '        �U�                    !       &        T&       '        �T�                    !       &        Q&       '        �Q�                    !       &        R&       '        �R�                                    U        !        �U�                                	        U	               S               U               �U�                          f        0�f       f        1�                                   P       h        V                      M       R        PR       V        TV       a        \                      ~      �       U�      �       \�              �U�                 ~      �       0�                  �      �       P                   ?      F       0�F      Y       V                  a      f       p } �                    �      �       U�      �       �U�                      �      �       U�      �       S�      �       �U�                        �      �       S�      �       �U $ &( �i     "��      �       S�      �       �U $ &( �i     "�                          �       U�      �       �U�                          �       T�      �       �l                        �             U             T      ~       ]~             �U�                      �      �       T�      |       \|             �T�                       )      +       V4      K       Vt      z       Vz             P                        y       S                        ~      �       U�      �       T�      �       V�      �       �U�                      ~      �       T�      �       \�      �       �T�                    �      �       P�      �       T                  �      �       S                      U      g       Ug      r       Sr      ~       �U�                      /      9       U9      T       VT      U       �U�                      <      J       PJ      S       SS      U       P                    6       K        UK       x        S                             <       S<      Y       UY      Z       sX�Z      �       S                          ?       ^?      Z       ~�Z      �       ^                          O       ^        P^       h        ]h       n        Pn       �       ]�      �       P                  '      G       S                 V              ^                        �       �        P�       �        \>      B       PB      �       \                                     \       C       x�C      Y       tx�Y      Z       h�\      �       x�                    ~       �        V�       �        v��       �       V                V             V                   ^      j       Pj             S                      u      �       _�      �       ��             _                 �      �      	 p r (�                                      U       5        \5       6        �U�                                     
�       2        S2       6        P                                   0�       "        V                          �      �       U�      �       \�             U      .       \.      /       �U�                    �      �       S�      �       S                    �      �       p s ��      �       Q                    �             U      %       \                  �      %       S                        %       Q                   �      
       0�
      %       P                        �      �       U�      �       S�      �       v �      �       �T                      �      �       T�      �       V�      �       �T�                       �      �       uX��      �       sX��      �       v (��      �       �T(�                      y      �       U�      �       S�      �       �U�                      y      �       T�      �       V�      �       �UH                      y      �       Q�      �       \�      �       �Q�                      y      �       R�      �       ]�      �       �R�                     y      �       uX��      �       sX��      �       �U(�                        x       S                      V      s       Us             V             �U�                               S                      �      �       U�      S       VS      V       �U�                      �      �       T�      U       \U      V       �T�                  �      R       S                      D      W       UW      �       S�      �       �U�                      D      W       TW      �       V�      �       �T�                      W      �       U�      �       uX��      �       U                  n      �       \                          6      ;       U;      C       u 	��C      N       UN      =       \=      D       �U#	�#(�                      6      o       To      ?       ]?      D       ph                      6      o       Qo      C       _C      D       �Q�                    �      �       Q�      �       p                   l      A       ^                 h      ;       V                  �      �       P                          \      o       Vo      �       S�      �       V�      :       S:      D       pX�                       D       P                        �       �        U�       4       S4      5       v(�5      6       �U�                    �              V      3       P                   �              P      6       Q                   Z       i        Ri       �        p(                                   P       7        u(                                      U       "        S"       2        �U�                                    T       2        �T�                                        Q       +        V+       1        U1       2        �Q�                                        R       -        \-       1        Q1       2        �R�                                     U       "        S"       2        �U�                        2       :        U:       C        SC       G        UG       H        �U�                       2       :        U:       C        SC       G        UG       H        �U�                    H       T        UT       �        �U�                    }       �        P�       �        S                    X       Z        PZ       �        V                  $       D        �W                  $       D        R                    *       6        1�6       >        	��                       [       d        �Wd       k        p ��C     "k       m        q  $ &��C     "m       o        0�                          �       U�      �       �U�                      4      K       UK      N       SN      }       �U�                    4      R       TR      }       �T�                    4      R       QR      }       �Q�                   S      b       0�b      }       P                     S      b       ����b      h       Tj      }       T                   S      b       0�b      }       R                 b      b       0���b      b      
 0��0���b      }       0��0��0��                    �      �       U�      �       u}�      4       U                     �      �       0��      �       Q�             q�      4       Q                    �      �       U�      �       �U�                <      <       ȟ                  7      �       \                �      <      ) D,f     �ԓe     ��P,f     �4%�                  <      <       P<      �       S                 <      �       ^                 <      �       V                      D      [       _[      ~       �~      �       _                    '      =       P>      S       P                            a       �        U�              S             u x "�             u x "#�             u x "�             S      ,       U                       a       j        Tj       q        t z "�      !       t z "#�!      ,       t z "�                     a       j        0�j              Z      !       z�!      ,       Z                    �              X             x�             X                   �       �        0��       ,       Y                    �       �        s 2$@(f     "�p�p���       �       2 s 2$@(f     "�s 2$A(f     "�s 2$B(f     "��                    �       �        Y�       ,       P                   �       �        p��8X,f     �&��       �       " s 2$B(f     "��8X,f     �&�                   �       �        p��8`,f     �&��       �       " s 2$A(f     "��8`,f     �&�                 �       �       " s 2$@(f     "��8h,f     �&�                                      U       ^        U`       a        U                                       T       )        t y "�)       [        t y "1�`       a        t y "�                                     0�       )        Y`       a        Y                 [       `        0�                        1       7        z 2$@(f     "�r�r��7       :        z 2$@(f     "�R�P��:       =       % z 2$@(f     "�z 2$A(f     "�P��=       [       2 z 2$@(f     "�z 2$A(f     "�z 2$B(f     "��                   1       7        r�3%�;$�7       [        z 2$B(f     "�3%�;$�                   1       7        r�2%�5$�7       [        z 2$A(f     "�2%�5$�                   1       V        z 2$@(f     "�3%��V       `        R                 @     @      1�                 @     @      
���                        �0B     1B      U1B     	1B      T	1B     1B      �U�1B     1B      U                  �0B     �0B      P                    �0B     �0B      U�0B     �0B      �U�                      /B     \/B      U\/B     �/B      S�/B     �/B      �U�                                                  /B     6/B      T6/B     `/B      P`/B     c/B      �T�c/B     h/B      Ph/B     j/B      Tj/B     o/B      Po/B     q/B      Tq/B     v/B      Pv/B     x/B      Tx/B     }/B      P}/B     /B      T/B     �/B      P�/B     �/B      T�/B     �/B      P�/B     �/B      T�/B     �/B      P�/B     �/B      �T�                 �/B     �/B      P                 �/B     �/B      s 8$p �!�                                              /B     6/B      T6/B     `/B      P`/B     a/B      �T�a/B     h/B      Ph/B     j/B      Tj/B     o/B      Po/B     q/B      Tq/B     v/B      Pv/B     x/B      Tx/B     }/B      P}/B     /B      T/B     �/B      P�/B     �/B      T�/B     �/B      P�/B     �/B      T�/B     �/B      P                                �@     @                     �       �       �                             �      �      �      �                      E      E      H      �                      �      �      �      �                      �      �      �      �                      �      �      �      �                      @      �      �      ]                      �      �      �      �                      �      �      �      �                             �      �      S                      �                  9      ;      G                      �      L	      M	      U	      V	      X	      Y	      ^	                      �      �      �      L	      M	      U	      V	      X	      Y	      ^	                      �	      �	      �	      �	      �	      �	      �	      �	                      o            T      �                                    5       �                       �       �       �       Z      _      h                      �      6      =      A                      F      �      �                                        �      �      �      $                            p      q      }                      �
      �
      �
      �
      �
      �
                      �Z@     �Z@     �Z@     �[@                     �Z@     [@     [@     )[@     G[@     �[@                     ]d@     bd@     ed@     4e@                     Df@     �f@     �f@     �f@     �f@     �f@     �f@     �f@     �f@     �f@                     	n@     mn@     nn@     sn@                     �W@     �y@                                                 )       1                                         #      '      +      .      <      ?      E                      '      +      .      <      C      E                      �      �      �      �      �      �                      �      �      �      �      �      �                      �      �      �      �                      �       �       �       �                                     I       p       r                              �       �       �       �       �       :                      n      q      �      5                      �      �      �      �                      �      �      -      /      3      �                      �      �      �      �            �      �                            2      2      4      ;      C      ~	      	      �	                      �	      �	      �	      �	      �	      B      C      H                      x      �      �      �      �                             �      �      �                            H      V      X      f      h      �      �      T      U      Z                      X      f      h      y      ~      �      �      H                      �      �      �      �      �      �      �      �      �      R      S      X                      �      �      �      �      �      �      �      �      �      �      �      ?                      �      �      �      �      �      �      �      �      �      �      �      �      �      �                      �      �      �      �      �      �      �      �      �      �      �      �                      �      �      �      �      �      �      �                  �      �      �                      �      �      �      �      �                              �                      �      �      �      �      �      �      �      �      �      �                      �                                        )      V      W      d                      �      �      �                  M                                                                  2       2       3       :                       �      �      �      5                      ��@     ��@     ǝ@     �@     ��@     ��@                     �@     �@     �@     �@     �@     �@                     &�@     &�@     '�@     I�@                     b�@     l�@     p�@     p�@                     ��@     ��@     ��@     ��@                     Ο@     Ο@     ϟ@     �@     �@     �@                     �@     �@     �@     .�@     3�@     @�@     G�@     J�@                     ��@     ��@     ��@     ��@     ¥@     ǥ@                     #�@     '�@     V�@     �@                     �@     ��@                           <      =      C                      4      4      :      S                             i       j       �       �       �                       Z      e      o      o      p      �      �                                         @      @      G      N                      A      H      N      �      �      �                      n      n      p      Z      [      ^      `      f                      J      �      �      �                      �       �       �       �       �       �       �                   )                      U      _      j      w                      |      �      �      �                      �      �      �      �      �      �      �      �                      �       �       �       �                       �      �      �      �      �                            G	      G	      J	      �	                      y      �      �      ,      .      4                      I      �      �      �      �      �                      ^      ^      f      H      P      Q                      �      �      �      �                      �      �      �                             �       �       �       �                       �       �       �       �       �       �                       �      �                                  �      �      �      G                      �      �      �      $                      �      �      �      �                      |      �	      �	      �	                      |      |      ~      �                                  R      �                      f      i      l      &                      *      -      0      �      �      �                      �      �      �                            I      L      O      �                      �      �      �      <      A      D                      �      �      �      �      �      �                      �      �      �      3      ;      >                      V      Y      \      �      �      �                      y       �       �       �       �       �                       �      �      �      o                                    $       )       _       g                       i
      i
      k
      �
                      �      �      �      �                      Z      ]      b      �      �      �      �                                                 !       $       )       *       /       0       ?       E       K                             #      )      8      <      B                      �      �      �      �      �      �                      :       D       O       �       �       �                       G      O      V      r      u                                                    $       $       &       D                       H       O       [       [       [       o                       /B     /B     /B     �/B                     /B     1B     @     @                     �BB     !CB     #CB     ,CB                     DB     �DB     �DB     �DB                     �>B     �DB     �DB     �DB     �DB     vEB     vEB     �EB     �EB     �EB     �EB     �EB     �EB     �EB      FB     �FB     �FB     �FB     �FB     �FB     �FB     �GB     �GB     �HB                             �  �  	  '	  7	  	P	  `	  
>7  4  �	  �	  ��  M6  �#  @  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �      .%   �4   #'   
   �5       h   �&   =   �
   �   3*      +7   �%   �:   �   �!   �    �   ,   �%   ?2   ?   Z$   w&   �   �   x5   >>   m      K,   >	   �(   O3   e   �<   B   �%   �   	+   o   �   MB   �0   n   �   �7   V2   �    e1   R   �   �      �	   �   �   �   �9   �'   �<   J&   �   �0   �4   	   ?A      $   �5      S   T
   �+   �   �.   �   4   �	   1   �&   �   t:   #&   s2   O4   z6   �   �   6-   �@   �5   �   0   �8   I/   ;   ;    1(   �+   U   �%   	*   v*   ^   q       �6   �   �   G   "
   /$   1   
A   �0   �8      �;   +   �   �&   �   F*   �?   5&   )#   F   �-   	C   ;   Y   t   �2   B   �C   �   �)   �!   �   4    0   �   2   (   �   t;   �   �   04   K   ?   (   7   �   �,   �   �7   :;   1   C   �$   p   \   �   *      k%   �=   �       J!   �A   �   �	   �;   �   '   �   -   j   �   pA   �C   `4   �    e	   5'      �      �0   w   �   L   �	      �@   �   �   �A   .   Z)   =
   �   ^   SC   �
   t<   �      T      P"   �   d3   r@   �   k   Y    �   �   B   �(   �   O   �@   �   j   �1   W>   �B   x   �.   �    Q    0   /   �   �?      �   �#         �   ^   �=   �3   �         �   !   �:   e   c-   J   eB      �/   �$   5)   z7   0   �   O   �   m$   iC   �   �.   �A   -   �   `/   �      :+   �/   Z?   H-   �<   �?   �%   �=   �   )   g      �!   �=   y   ;5   ,   �:   ~   3    �6   �   x4   >$   1B   �   �(   �   �   @   H   V.   �   �=   5   �5   �   #   �6   !   �   �   >   9%   �8   �*   �2   �4   �*   �9   �   �#   -;   �!   �     �   '  f� v�    "  �"  �  C     ,+  �     ��Q  �`  ��     �  �*     ��"  ��  �}  ��>  �x  ��2  �+  �A  �=  �|  ��  �x  ��=  �"*  �y  ��  �P?  ��)  ��     "�)  '�3     �&  w9  =<  >A  ?P  AE  C_  E�  F5  GX1  I     3  �  �  �   W  "�  #�,  $�  %  (�  )�&  *�/  +>  -E  .:  /�  0S  2�  3�+  4$=  5P@  R�>  S  T�+  W<  X*  Y�  \    ]R+  ^  a�  b$6  c^(  �I:  ��  ��;  ��  �O7  ��3  ��  �$  ��9  �.  ��,  ��4  �  �t
  ��  ��>  �\8  �x  �F=  ��  ��#  �W0  ��1  ��  �>8  ��  �c   �"  �3     ;5  <�'  =�  >�B  Ae,  BA  C�  D�  K�  L.!  M�  N�%  P$1  Q�  R&  SO%  V�  W&?  X�  YZ  \�6  ]/9  ^/  _�"  a�  b�;  c�8  d�.  gk  h�-  i�2  j  m�
  n�
  o�1  p6<  ra  s8  tt  u�  xQ9  y�8  za.  {L  ~M  �7  �\6  ��   ��  �0@  ��2  �E  �[  �  �q  ��   ��  �%  ��     1/  �  	q'  
 9  ;/  w=  T  �%  i  �    >1  �B  �   �3  +   �  �  �5  _  �>   B  D  �  �    g
  !�  "�  #"  $�#  %fA  &N1  '�  (%  )�"  *�  +  ,3  -53  .Q  /�  0�6  1%  2D4  3  4{+  5g&  6J  7�*  8�'  9�,  :~  ;D%  <�.  =�  >�*  ?5  @�?  A�  B :  C]5  DJ)  E&  F�  G�<  H�7  IC3  J/  K�&  L�  M�0  N�$  O�,  P  Q�  R�  S8  T�'  U�+  V"  W�8  X�(  Y�,  Z�  \D?     �'    40  n5  m5  	Y  
�5  �  �  �2  "@  �(  �     <�(  ? +  @�9  Dj=  H�0  I2  J�  K\<  N�  R�!  `�0  a�0  b�  c�  g�  h (  i�?  j)A  m�?  q�B  uJ�  v�"  w^j  x�   {�,  |.,  ��  ��  �o5  ��6  ��  ��/  ��  �k  �n5  ��5  �m5  ��)  ��?  �   ��  �V*  ��  ��$     ^�'  _3  `�  d�-    �     �<  #w0  P	  `	  2�:  ?�  	�  	?
  �  �  G  T
%  "�'  
�I  s   �  �    �     �  ,�  -	  .'	  7	  /P	  `	  0>7  4  1�	  �	  �2�  3M6  �#  ˈ  �<  #4w0  2�:  ?5�  6	�  ?
  �  �  G  T7%  "8�'  7�9I  s   �  �  :�  ;�  <��     0  =@  
x�  >��  ??��  @�  	{�  �  &�  �  �    !��  AZ�  #�  '  2  B��  ��  !�  #�S   �  %3_  %�  'j�  �  x  ��  ��    &  (C3  B%�  &��  'D՘  (�l  *�  + 2�  �  �"�  $�z  #W�   %��  !+X{  1  "EiN  %&V  ((�r  ':�  f  ,)#�  Fw  #  .*#  2��  3�X  4�P  5��  6�a  7�  8��  9BF  :\v  ; �  <��  =��  >.�  ?�M  B��  C��  DSi  E�e  FF  G�Q  H&�  I�  J՛  K7�  L�F  M �  N`�  O�  Pr�  Q��  Rb�  S��  W�  Z��  ]��  `��  c�c  f+�  g*W  i	�  j߅  m¸  ��  �R ��  �R ��Y  �R ��Y  �R ���  ���  �fy     ��  Bc   �   �  $�     Ə  &R]  'x�  (:�  )N�  *��     ��  �O     �w  E�s     0�  ?�  ��  4�  U  �   �|  !۠  "�d  #e� $�  %��  &=�  '�W  (�p  )�  *��  +4�  ,i�  -�Q  ._i  /��  0�}  1v�  3�  4��  6PF  7Ew  9Iq  :i  ;�  =�f  A�y  B9�  C�i  D�}  FE�  G��  HV�  IΩ  J�j  Ko�  MI�  N��  O�U  P|�  Q�q  R�g  S�w  TZQ  U�q  Vd�  X�t  Y��  Z�o  [��  \��  ]u�  ^)�     D�  2�     "��  %��  *��  -K�  M�M  N>�  Oo�  R�     F�  �   @�  !�a     %�  �   �|     Y�  �n  �m     )�  *��  .��  ?��  @L�  AR�  B۟  CN�  E�H  F��  K�|  Mz  NՓ  O9�     ��  b��  e�  i_}  u��  x�  {��  ~��  ���  �h�  ���     rv  �_  m~   e�  $]�  &��     .,�  /��  0_�  1��  3�a     ��  ,e  -�`     tR  `�  %�  )��  -U|  gqn  k�H  ��j  ��e  ���  ���  ��  �y�  �jo  ��     ǔ  =�  >T  @w]  A|�  B��  C�  O1�     |`  ;�     ��  ��  ��  #F�  $�  %�i  &�R  'u  +��  0tH  2��  3T�  5D�  6Rs  7e�  :u�  \A�  ]Sj  `�w  ���  �'j  ��t  �>�  ��d  ��  �`F     �y  #={  ���  ��y  �~�  ��  �2�  �)H  ���  ���  ��j  �OV  �a\  ��K  �)�  ���  ��v  �	x     �|   ��  "�)  /��  0}K  1��  4��  6��  i�  l�3  o��  r�  u��     �H  "�     E�o  ��S     ��  �  :R  $��  %)�  &�  '.�  (X  )�K  *�  +�  ,��  . �  2�[  6��  :�|  ;�  <K�  =;�  ?��  A3�  Ba�  CFh  D��  E#�  F�Q  GC�  H�W  M��  N�v  Oҋ  P3�  Q�d  R9^  S �  T�c  V6�  WMe  X��  Y�G  Z��  [�\  ]�S  ^=�  _�J  `QW  a�i  b-�  c��  e��  f�  g�  hc  i��  jp�  k��  l��  m�n  oU�  pF�  q#`  ry�  s6y  tk�  us�  z~  {�  |�  }d�  ~5�  	�  ��  �C�  �l�  �$w  �B�  ���  ��M  �Az  �6�  ��  �V  ��g  �E�  ��X  ��l  ��  ��g  ���  �d�  �h�  ���  �Q_  ��`  ���  �B�  �|^  �X�  ��w  ���  �x�  ��_  �]c  �N�  � w  �׍  ��  ���  ���  ��x  ���  ���  �_�  ��x  ���  �P�  �Һ  �5�  ��r  ���  �ʲ  ���  ���  �+�  �Q�  �*}  �"�  �!�  ���  ���  ���  �P�  �	^  �dO  �Q�  �d�  �zG  �f  ���  �*�  ���  ���  �v  ��u  �y  ���  ���  �:�  �ʝ  �I�  ���  ��M  ���  �S�  ��R  �ܪ  �a�  ���  ��O  �ǫ  �w�  �!�  ���  �ۼ  ��  �v_  ���  �-V  �ԙ  ���  �_X  �'T  ���  ��  �b  ���  ��  �\l  ��S  �#D  �-Q  ��  ��b  �	�  �3�  �H�  ��b  ���  ��  ���  �ri  �-�  ��  ��c  �Y�  ��i  ���  ���  �7H  ��]  ���  ��t  ��  �`x  ��  �7�  �y�  �R  �5�  ���  �"�  ���  �w\  �d�  �.�  �wN  ���  ��`  ��  ��F  ��T  ��s  �2e  � �  �չ  ���  ���  ��\  �W�  �z�  ��  ���  �l  ��k  �ƌ  ���  �we  �M�  �f�  ��O  ��^  �ˁ  ���  ��  ��  ���  �Ӕ  ���  ��Y  ���  ��  �7�  �F�  �>D  ���  ���  �Ik  ���  �P�  ���  ��  �z�  �u�  ��H  �X�  �<L  ���  �[V  ���  �{F  �;O  ���  ���  �B�  ���  �n�  ��F  ��Y  ���  �*�  ��k  �+�  �^�  �MT  ���  ��z     +c  #�w     ��  ��  �  Q�    	     �  �  	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  �r  ��  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T %  "!�'   �"I  s   �  �  x�  #��  ?$��  %�  {�  �  %  
:�  &tR  	  '��  P%  "��  ��  ��    �%  $3_  �  &  !�S  f     b��  e�  i_}  u��  x�  {��  ~��  ���  �h�  ���     `�  %�  )��  -U|  gqn  k�H  ��j  ��e  ���  ���  ��  �y�  �jo  ��     #�  )�  *��  .��  ?��  @L�  AR�  B۟  CN�  E�H  F��  K�|  Mz  NՓ  O9�     ,e  -�`    �      #�  w  #    �      ��  P'  	  '	  7	  P	  `	  	`'  p'  	
��  �'  y��  �  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  $�     ;�  ��     ��  G�     ���  ���  ���  ���  � �  �.�  ��  ��  ���  �W�  ���  �u�  ���  ���  ���  ���  ��  ��     s�  ��   ��  #�    �#     3_  �  ��  x�  �  �  		  
'	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  ��  ?��  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  �  {�  �    v&     �  �  	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  ��  P'  `'  p'  	��  �'  y��   �  ��  ?��  !w+  "Ə  #�  A,  $@  5�  {�  �<  #w0  2�:  ?%�  &	�  ?
  �  �  G  T'%  "(�'  '�)I  s   �  �  c,  iN  *  +�  	@  
��  X{     �z  W�  !,0  :l�     �  ��  
�� `�  P�  ��  �  ��  �  ��  "o�  %��  ()�  +��  .�� 1=� 4-� 7�� :3�  =� @��  C��  F��  I�  L.�  O��  R�� Ur�  XC�  [��  ^z�  a��  d��     &R]  'x�  (:�  )N�  *��     ^�  �  r�   A�    P.     ��  P'  	  '	  7	  P	  `	  `'  p'  	��  �'  y��  ��  ?��   �  �  �<  #!w0  2�:  ?"�  #	�  ?
  �  �  G  T$%  "%�'  $�&I  s   �  �  :�  
tR  �  '�  (>7  4  )�	  �	  �*�  +M6  �#    	��  P%  iN  �  �   @  !  # $,) %��  &-��  '.�  (S�  )4   �7     D�  �  E�  F	  G'	  7	  HP	  `	  I>7  4  J�	  �	  �K�  LM6  �#  7��  MP'  N`'  p'  	O��  �'  yP��  8��  ?Q��  Rw+  ˈ  �<  #?w0  2�:  ?S�  T	�  ?
  �  �  G  TU%  "V�'  U�WI  s   �  �  X�  Y�  ��     
x�  <�  	{�  �  �r  �  :�  tR    P%  "��  ��  ��    �%  $3_  �  &  !�S  f  !#�  Zw  #  #K � %9�2  '0  (:c )�z  W�  *� + �H  [j�  "�  -B� !�  ."�	 0#@  1$��  2%��  3;X{  J  4&� 5'�2  7@� 8=�2  9(iN  ;)�  =*| ?+E3  @A� A-&�  ,�    B.#  C/ D\ 
 E]��  G>� H^Z�  _��  �3  0x  _%1�  &2��  '`՘  (3�l  *4�  +52�  Ia�
 K6�    5�  ^�  �  r�   A�     7     � � !( $; '� (� +� 0m 2{ 5y 7 9 <� =M	     � � � !� #A $l %m &� (�    ��  .,�  /��  0_�  1��  3�a    �K     �<  #w0  P	  `	  2�:  ?�  		�  
?
  �  �  G  T%  "�'  �I  s   �  �  {�    �N     "��  #P'  $	  %'	  7	  &P	  `	  '`'  p'  	(��  �'  y)��  *�  	� x�  �  +�  ,>7  4  -�	  �	  �.�  /M6  �#  0��  ?1��  �<  #2w0  2�:  ?3�  4	�  ?
  �  �  G  T5%  "6�'  5�7I  s   �  �  8�  {�  �  
@  � 9�  !X{  -  :iN    �  | !�r  �  :�  tR  ��  P%  "��  ��  ��    �%  $3_  �  &  !�S  f  " $ #�z  W�  %ˈ  ;�       JV     �  &�  '	  ('	  7	  )P	  `	  *>7  4  +�	  �	  �,�  -M6  �#  %�  ˈ  �<  #.w0  2�:  ?/�  0	�  ?
  �  �  G  T1%  "2�'  1�3I  s   �  �  4�  5�  6��     7iN    	�  8�9  
0  �H  j�  "�  �z  {�  W�  � �S  #�  '  2  �   ��  x�  9��  ?:��  ;�  �  %  %3_  K � !� "#�  <w  #  %!�r  :�  =3  "��  ��     f  &#x  >��  ��  %"�  �  #98 :� �$E3      /� 0] 2�   {b     ��  	  '	  7	  P	  `	  ?��  �w  �  �  >7  4  �	  �	  ��  M6  �#  E�s  rv  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  _;  	�H  j�  "�  
 �	    �_  m~   e�  $]�  &��    �i     ?��  @	  A'	  7	  BP	  `	  ?C��  7��  DP'  E`'  p'  	F��  �'  yG��  H�?  x�  �  I�  J>7  4  K�	  �	  �L�  MM6  �#  �<  #Nw0  2�:  ?O�  P	�  ?
  �  �  G  TQ%  "R�'  Q�SI  s   �  �  4�  {�  �  T@  �r  	�  :�  UtR  
  V��  P%  "��  ��  ��    �%  $3_  �  &  !�S  f  ˈ  W�  X�     Y�@  0   :� �  !@  "��  #6X{  K  $� %8 &5iN  (�  *>� +�2  ,=� .� 0<� 1E3  2!&�   �    3"#  4;�
 7#�H  Zj�  "�  9%�z  $W�  ;,��  [Z�  9��  �3  &x  9%'�  &(��  '\՘  ()�l  **�  ++2�  �  �-�  =0� /K .� @1#�  ]w  #  E2�A  I3| LX1 ��  �  �I1 �$% �L  ��! �* ��(     �- � � 	Z! 
�$ ;* ) �# � K.   " H" � U/ i"  . !�" "�. #0% '1 (�' )�/ /�$ 0�) 1�' 2x, 3�" 9�+ ?n* @�# AI# B�, E�  H�( [�* `7 av- b{% c<) d�0    k/  & �, $ �! � ` �/ 9$  g !�0 "}  #�0 $@ %�, &s ?o$ @/ A�% B�! CM& D�& EH( F90 Gi. HA+ I� JF, K* L�) M�' N(     �& �    .�     �  x�  �  �  	   '	  7	  !P	  `	  ">7  4  #�	  �	  �$�  %M6  �#  &��  ?'��  �<  #(w0  2�:  ?)�  *	�  ?
  �  �  G  T+%  ",�'  +�-I  s   �  �  .�  /{�  �  0@  	�H  j�  "�  1�9  h2 ��  
  !�  #�S  �%   �  %3_  %�  �  (D  2Z�  3��  x  ��  ��    &  (4tR  5��  P%  3%�  &��  '6՘  (�l  *�  +2�   x3    M2 Y3 �3   l�     %�  x�  �  &�  '	  ('	  7	  )P	  `	  *>7  4  +�	  �	  �,�  -M6  �#  .��  ?/��  �<  #0w0  2�:  ?1�  2	�  ?
  �  �  G  T3%  "4�'  3�5I  s   �  �  6�  {�  �  7@  	0  
ˈ  8�  9�  :��     ;�9  �   �  YG  h2 ��    !�  #�S  �%   �  %3_  'j�  �  (D   ��  !$X{  +  "�z  W�  $� K � &"�r  :�  <tR    P%  "��   ��  !  f  )##�  =w  #  /�3 0T6 1�5 2~5 3a4 4�3 5)6 6�4 86 9B6 :4 ;4 <�6 ��4    � � � !� #A $l %m &� (�   ��     �  �  	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  ��  P'  `'  p'  	��  �'  y��  K � �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  � I  s   �  �    
3_  	�  �S  �%   !��  "x�  #��  ?$��  %�  &{�  �  %    l�     �  �  	  '	  7	  P	  `	  	>7  4  
�	  �	  ��  M6  �#  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  qJ     �6 �6 �7 �7 �7 17 C7 �6   ?�     �  �  		  
'	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  ��  ?��  w+  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  �  '8 38   �     ��  P'  	  	'	  7	  
P	  `	  `'  p'  	��  �'  y��  �  �  >7  4  �	  �	  ��  M6  �#  ��  ?��  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  �  �2   iN  !   ��  !X{    &9   ǫ     �  �  	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  ��  P'  `'  p'  	��  �'  y��  ��  ?��  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  �  @  	0  ��< �	y= �	�< �
5=   ��     �  �  	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  ��  P'  `'  p'  	��  �'  y��  w+  �  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �   � !�  "	@  #
��    {�     ��  P'  	  '	  7	  P	  `	  `'  p'  	��  �'  y��  �  �  >7  4  �	  �	  ��  M6  �#  ��  ? ��    
C ?
  !�J 	"�D #*F �R  %$w+  '%Ə  &�  A,  (	�<  #w0  2�:  ?'�  (	fT  �  G  T)%  "*�'  )�+I  s   �  �  )
@  *��  +X{  ,,�2  -� .-�  /�  1iN  .  /�  3�z  0{�  W�  410  :)G ;�B ��A ��E    !J KI �G J }C LJ D �C �A  $C !�H "�A #�A $�D &�J 'NG (�G )-D *�J +;B ,#A -YA .�B /IC 0�G 1�I 2H 3[E 4UD 5�F 6�B 7�C 8�E 9�D :�C ;�D <OF =�B >�H ?}H @tI A�I B�F C3H DfJ EI F�H G�G K�E LBI MD N�E RAE S�A T	F U�I XyD YsF ZcI [qB \�H ]bB _�I `B a+B    �  ;5  <�'  =�  >�B  Ae,  BA  C�  D�  K�  L.!  M�  N�%  P$1  Q�  R&  SO%  V�  W&?  X�  YZ  \�6  ]/9  ^/  _�"  a�  b�;  c�8  d�.  gk  h�-  i�2  j  m�
  n�
  o�1  p6<  ra  s8  tt  u�  xQ9  y�8  za.  {L  ~M  �7  �\6  ��   ��  �0@  ��2  �E  �[  �  �q  ��   ��  �%  ��    ��     �  �<  #w0  P	  	`	  2�:  ?
�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  �V  �V     eK 5K  K    �|   ��  "�)  '�3  /��  0}K  1��  4��  6��  i�  l�3  o��  r�  u��    '�     �  �  	  	'	  7	  
P	  `	  >7  4  �	  �	  ��  M6  �#  ��  P'  `'  p'  	��  �'  y��  ��  ?��  �K 0    ��     �  �  	�  
	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  ��  P'  `'  p'  	��  �'  y��  ��  ?��  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  iN     �  !X{    @  I�L   f�     M %  "�'  �I  s   �      ��     ��  	  '	  7	  P	  `	  ?	��  �<  #
w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  �    t�     �  �  	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  	��  P'  `'  p'  	��  �'  y��  ��  ?��  �  LQ �\  oO w+  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T %  "!�'   �"I  s   �  �  #@  $�   
iN  %  &�  !@  "X{    $'0  _|N b�N d�P feR h/T jS    DQ 5U U fO DP 	�O 
�Q �Q �T �S �Q 1R �N qN �M �S nU lM �U �N bQ /Q �S �M �T &P R OM  �M !�R "�U #�U $�O %P &�O '�U (�R )U *�Q +�T ,1O -Q .CM /�P 0@O 1�M 2�O 3�Q 4�U 5T 6VQ 7�O 8�P 9�R :�M ;�O <�U =4N ><U ?IN @8P A[O B�N CLO DT E�Q F�S G`M H�S I�S J�S K�O L�S M%R N Q ON P[U Q<R R�P S�Q T�O   ��     �  �  	  '	  7	  	P	  `	  
>7  4  �	  �	  ��  M6  �#  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  @  ��  X{      ��     ��  P'  	  '	  	7	  
P	  	`	  `'  	p'  	��  �'  y��  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  iN    �      ��     5��  6P'  7	  8'	  7	  9P	  `	  :`'  p'  	;��  �'  y<��  2�  x�  �  =�  >>7  4  ?�	  �	  �@�  AM6  �#  3��  ?B��  �<  #Cw0  2�:  ?D�  E	�  ?
  �  �  G  TF%  "G�'  F�HI  s   �  �  1�  {�  �  I@  	#�  Jw  #  
� ˈ  K�  L�  M��      N�9  !0iN    �  #�  $/X{  ?  %�H  j�  "�  &�z  W�  '0  )OZ�  #�  '  2  P��  ��  !�  #�S   �  %3_  �  x  ��  ��    (Q3  P%�  & ��  'R՘  (!�l  *"�  +#2�  ,$E3  .%| 0&@  1'��  2(�2  4+� *K )� 6-�r  ,:�  f  ;.� x�W yI[   �    �  �  	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  ��  P'  `'  p'  	��  �'  y ��  ��  ?��  �  LQ !�\  oO #b " ^ #�] $�J %�D &�] '�a 	(�a 
)Na *�] +�] ,�] -�a |g  
h  $.B^ 	/�` 0*F 1Q` 2.^ 3P^ '	�<  #w0  2�:  ?4�  5	�  ?
  �  �  G  T6%  "7�'  6�8I  s   �  �  )9Ə  :�  A,  +;�9  ,iN  <  =�  -
�  .>X{    /�H  ?j�  "�  0�z  @{�  W�  10     �` A` �] 3a �a �a �_ �_ �^ sa �^ �^ 5` �^ _  �] !�^ "|^ #�] $Ca %` &�_ '^    �a a �` 	�^ 
�_ -_ T_ \] d^ n`   �      x    �w  �  #�  $	  %'	  7	  &P	  `	  '>7  4  (�	  �	  �)�  *M6  �#  E�s  	x�  +��  ?,��  �<  #-w0  2�:  ?.�  /	�  ?
  �  �  G  T0%  "1�'  0�2I  s   �  �  3�  {�  �  ��  4Z�  #�  '
  2  5��  ��  !�  #�S   �  %3_  %�  '6j�  �  x  ��  ��    &  (7tR  8��  P%  5%�  &��  '9՘  (�l  *�  +2�  �  ��   � K � "�r  !:�  f    !    �w  �  &�  '	  ('	  7	  )P	  `	  *>7  4  +�	  �	  �,�  -M6  �#  E�s  	x�  .��  ?/��  �<  #0w0  2�:  ?1�  2	�  ?
  �  �  G  T3%  "4�'  3�5I  s   �  �  6�  {�  �  
ˈ  7�  8�  9��     ��  :Z�  #�  '  2  ;��  ��  !�  #�S   �  %3_  %�  '<j�  �  x  ��  ��    &  (=3  ;%�  &��  '>՘  (�l  *�  +2�  �  ��  !�  K � #�r  ":�  f  !$#�  ?w  #    k+    �  %�  &	  ''	  7	  (P	  `	  )>7  4  *�	  �	  �+�  ,M6  �#  -��  .P'  /`'  p'  	0��  �'  y1��  # �<  #2w0  2�:  ?3�  4	�  ?
  �  �  G  T5%  "6�'  5�7I  s   �  �  $iN    8�  	x�  9��  ?:��  ;�  {�  �  ��  <Z�  #�  '
  2  =��  ��  !�  #�S   �  %3_  %�  '>j�  �  x  ��  ��    (?tR  @��  P%  =%�  &��  'A՘  (�l  *�  +2�  �  ��  � K �   | #"�r  !:�  f  �
�j ��f   �J    �w  �  #�  $	  %'	  7	  &P	  `	  '>7  4  (�	  �	  �)�  *M6  �#  E�s  	x�  +��  ?,��  �<  #-w0  2�:  ?.�  /	�  ?
  �  �  G  T0%  "1�'  0�2I  s   �  �  3�  {�  �  ��  4Z�  #�  '
  2  5��  ��  !�  #�S   �  %3_  %�  '6j�  �  x  ��  ��    &  (7tR  8��  P%  5%�  &��  '9՘  (�l  *�  +2�  �  ��   � K � "�r  !:�  f    �U    x�  �  (�  )	  *'	  7	  +P	  `	  ,>7  4  -�	  �	  �.�  /M6  �#  0��  ?1��  �<  #2w0  2�:  ?3�  4	�  ?
  �  �  G  T5%  "6�'  5�7I  s   �  �  8�  {�  �  	#�  9w  #  K 
� ˈ  :�  ;�  <��     =�@  �r  �  :�  >tR    P%  "��  ��  ��    �%  $3_  �  &  !�S  f  &  'iN  ?�  "��  �  lv  $#��  @Z�  A��  ��  %�  'Bj�  �  x  A%�  &��  'C՘  ( �l  *!�  +"2�  �  �$�  &%� (D�l +Km    ��  �  Q�    Pf    �w  �  �  	   '	  7	  !P	  `	  ">7  4  #�	  �	  �$�  %M6  �#  E�s   �<  #&w0  2�:  ?'�  (	�  ?
  �  �  G  T)%  "*�'  )�+I  s   �  �  x�  ,��  ?-��  .�  /{�  �  ��  0Z�  
#�  '	  2  1��  ��  !�  #�S   �  %3_  %�  '2j�  �  x  ��  ��    &  (3tR  4��  P%  1%�  &��  '5՘  (�l  *�  +2�  �  ��    �n    �  '�  (	  )'	  7	  *P	  `	  +>7  4  ,�	  �	  �-�  .M6  �#  /��  0P'  1`'  p'  	2��  �'  y3��  4k/ 5�  |  M 6%  "7�'  6�8I  s   �    % �<  #9w0  2�:  ?:�  ;	�  ?
  �  �  G  T6�  $iN  	  <�  x�  =��  ?>��  ?�  
{�  �  @  &X{  ,   ��  @Z�  �%  A��  ��  !�  #�S   �  %3_  %�  'Bj�  �  x  ��  ��    (CtR  D��  P%  A%�  &��  'E՘  (�l  *�  +2�  �  ��  "!�  K � %#�r  ":�  f  2p     & �, $ �! � ` �/ 9$  g !�0 "}  #�0 $@ %�, &s ?o$ @/ A�% B�! CM& D�& EH( F90 Gi. HA+ I� JF, K* L�) M�' N(   o�     ��  !P'  "	  #'	  7	  $P	  `	  %`'  p'  	&��  �'  y'��  M (%  ")�'  (�*I  s   �    
x�  �  +�  ,>7  4  -�	  �	  �.�  /M6  �#  0��  ?1��  �<  #2w0  2�:  ?3�  4	�  ?
  �  �  G  T(�  5�  	{�  �  �r  �  :�  6tR    7��  P%  "��  ��  ��  �%  $3_  �  &  !�S  f   ��  8Z�  9��  ��  %�  ':j�  �  x  9%�  &��  ';՘  (�l  *�  +2�  �  ��    ��    �  (�  )	  *'	  7	  +P	  `	  ,>7  4  -�	  �	  �.�  /M6  �#  'iN    �<  #0w0  2�:  ?1�  2	�  ?
  �  �  G  T3%  "4�'  3�5I  s   �  �  6�  0  & 
x�  7��  ?8��  9�  	{�  �  ��  :Z�  #�  '  2  ;��  ��  !�  #�S   �  %3_  %�  '<j�  �  x  ��  ��    (=tR  >��  P%  ;%�  &��  '?՘  (�l  *�  +2�  �  ��  K � !&�   �    "E3   #� "%�r  $:�  f  iAt j�s   	�    �  %�  &	  ''	  7	  (P	  `	  )>7  4  *�	  �	  �+�  ,M6  �#  #iN    �<  #-w0  2�:  ?.�  /	�  ?
  �  �  G  T0%  "1�'  0�2I  s   �  �  3�  0  $ 
x�  4��  ?5��  6�  	{�  �  ��  7Z�  #�  '  2  8��  ��  !�  #�S   �  %3_  %�  '9j�  �  x  ��  ��    (:tR  ;��  P%  8%�  &��  '<՘  (�l  *�  +2�  �  ��   � K � "�r  !:�  f    ?�    x�  �  $�  %	  &'	  7	  'P	  `	  (>7  4  )�	  �	  �*�  +M6  �#  ,��  ?-��  �<  #.w0  2�:  ?/�  0	�  ?
  �  �  G  T1%  "2�'  1�3I  s   �  �  4�  {�  �  	�  5k/ 6�  |  # ��  7Z�  #�  '
  2  8��  ��  !�  #�S   �  %3_  %�  '9j�  �  x  ��  ��    &  (:tR  ;��  P%  8%�  &��  '<՘  (�l  *�  +2�  �  ��   � K � "�r  !:�  f  &qv '�v )�u *ou   ռ    �  )�  *	  +'	  7	  ,P	  `	  ->7  4  .�	  �	  �/�  0M6  �#  '��  1P'  2`'  p'  	3��  �'  y4��  #�  5w  #  ˈ  �<  #6w0  2�:  ?7�  8	�  ?
  �  �  G  T9%  ":�'  9�;I  s   �  �  <�  =�  >��     $iN  	  ?�  
0  ��  @Z�  #�  '  2  x�  &��  ?A��  B�  {�  �  C��  ��  !�  #�S   �  %3_  %�  'Dj�  �  x  ��  ��    (E3  C%�  &��  'F՘  (�l  *�  +2�  �  ��   �2  "�r  !:�  f   #| !%X{  .  $hw %* �qy ��z ��y ��w   k�    +�?  �w  �  ,�  -	  .'	  7	  /P	  `	  0>7  4  1�	  �	  �2�  3M6  �#  E�s  ˈ  �<  #4w0  2�:  ?5�  6	�  ?
  �  �  G  T7%  "8�'  7�9I  s   �  �  :�  ;�  <��     =�9  	@  M 7
  | x�  >��  ??��  @�  {�  �  A�    !*iN  "�z  W�  %"��  BZ�  �%  )��  ��  !�  #�S   �  %3_  %�  'Cj�  �  x  ��  ��    (D3  )%�  &��  'E՘  (�l  * �  +!2�  �  �#�  '&� %K $� )(�r  ':�  f  i�{   ��    x�  �  �  	  '	  7	   P	  `	  !>7  4  "�	  �	  �#�  $M6  �#  %��  ?&��  �<  #'w0  2�:  ?(�  )	�  ?
  �  �  G  T*%  "+�'  *�,I  s   �  �  -�  .{�  �  iN    /�  ��  0Z�  
#�  '	  2  1��  ��  !�  #�S   �  %3_  %�  '2j�  �  x  ��  ��    (3tR  4��  P%  1%�  &��  '5՘  (�l  *�  +2�  �  ��    ��    -��  .P'  /	  0'	  7	  1P	  `	  2`'  p'  	3��  �'  y4��  x�  �  5�  6>7  4  7�	  �	  �8�  9M6  �#  :��  ?;��  �<  #<w0  2�:  ?=�  >	�  ?
  �  �  G  T?%  "@�'  ?�AI  s   �  �  B�  {�  �  �r  	�  :�  CtR  
  D��  P%  "��  ��  ��    �%  $3_  �  &  !�S  f  ˈ  E�  F�     (iN  G�  0   @  !)X{  7  "* #�z  W�  %HZ�  +��  ��  %�  'Ij�  �  x  +%�  &��  'J՘  (�l  * �  +!2�  &"�  �#�  ($| *'� &K %� N �� �� �	@~ �	�~    ��  ��  ��  ��  #F�  $�  %�i  &�R  'u  +��  0tH  2��  3T�  5D�  6Rs  7e�  :u�  \A�  ]Sj  `�w  ���  �'j  ��t  �>�  ��d  ��  �`F    �    �  &�  '	  ('	  7	  )P	  `	  *>7  4  +�	  �	  �,�  -M6  �#  %iN    �<  #.w0  2�:  ?/�  0	�  ?
  �  �  G  T1%  "2�'  1�3I  s   �  �  4�  ˈ  5�  6�  7��     
x�  8��  ?9��  :�  	{�  �  ��  ;Z�  #�  '  2  $��  ��  !�  #�S   �  %3_  %�  '<j�  �  x  ��  ��    (=3  $%�  &��  '>՘  (�l  *�  +2�  �  ��  | !�  K � ##�r  ":�  f    �    x�  �  "�  #	  $'	  7	  %P	  `	  &>7  4  '�	  �	  �(�  )M6  �#  *��  ?+��  �<  #,w0  2�:  ?-�  .	�  ?
  �  �  G  T/%  "0�'  /�1I  s   �  �  2�  {�  �  �r  	�  :�  3tR  
  4��  P%  "��  ��  ��    �%  $3_  �  &  !�S  f  � K �  ��  5Z�  6��  ��  %�  '7j�  �  x  6%�  &��  '8՘  (�l  *�  +2�  �  �!�    $    �w  �   �  !	  "'	  7	  #P	  `	  $>7  4  %�	  �	  �&�  'M6  �#  E�s  ��  (Z�  #�  %�<  #)w0  2�:  ?*�  +	�  ?
  �  �  G  T,%  "-�'  ,�.I  s   �  �  '  2  
x�  /��  ?0��  1�  	{�  �  2��  ��  !�  #�S   �  %3_  %�  '3j�  �  x  ��  ��    &  (4tR  5��  P%  2%�  &��  '6՘  (�l  *�  +2�  �  ��  �r  :�  f    I    x�  �   �  !	  "'	  7	  #P	  `	  $>7  4  %�	  �	  �&�  'M6  �#  (��  ?)��  �<  #*w0  2�:  ?+�  ,	�  ?
  �  �  G  T-%  ".�'  -�/I  s   �  �  0�  {�  �  	�  ��  1Z�  #�  '
  2  2��  ��  !�  #�S   �  %3_  %�  '3j�  �  x  ��  ��    &  (4tR  5��  P%  2%�  &��  '6՘  (�l  *�  +2�  �  ��  �r  :�  f  "1� *�� �ۀ   �    x�  �  �  	  '	  7	   P	  `	  !>7  4  "�	  �	  �#�  $M6  �#  %��  ?&��  �<  #'w0  2�:  ?(�  )	�  ?
  �  �  G  T*%  "+�'  *�,I  s   �  �  -�  {�  �  
M *	  iN    .�  ǔ  ��  ��  ��  �%  $3_  �  &  !�S   �  (/tR  0��  P%  1��  ��  %�  '2j�  �  x  1p�  �l  �  !�r  :�  f  Q��    =�  >T  @w]  A|�  B��  C�  O1�    6(    �  )�  *	  +'	  7	  ,P	  `	  ->7  4  .�	  �	  �/�  0M6  �#  ˈ  �<  #'w0  2�:  ?1�  2	�  ?
  �  �  G  T3%  "4�'  3�5I  s   �  �  6�  7�  8��     9�9  %iN    :�  	0  �z  
{�  W�  x�  ;��  ?<��  =�  �  &X{  .   >Z�  #�  '  2  ?��  ��  !�  #�S   �  %3_  %�  'j�  �  x  ��  ��    (@3  ?%�  &��  'A՘  (�l  *�  +2�  ! �  �!�  ##�r  ":�  f  $$�A    �9    x�  �  $�  %	  &'	  7	  'P	  `	  (>7  4  )�	  �	  �*�  +M6  �#  ,��  ?-��  �<  #.w0  2�:  ?/�  0	�  ?
  �  �  G  T1%  "2�'  1�3I  s   �  �  4�  {�  �  	ˈ  5�  6�  7��     #iN  
  8�  0  �z  W�  9Z�  #�  '  2  :��  ��  !�  #�S   �  %3_  %�  'j�  �  x  ��  ��    (;3  :%�  &��  '<՘  (�l  *�  +2�  " V  %"�r  !:�  f  )�� *5� -�� ��� �Ӆ   II     ��  !P'  "	  #'	  7	  $P	  `	  %`'  p'  	&��  �'  y'��  (�?  x�  �  )�  *>7  4  +�	  �	  �,�  -M6  �#  .��  ?/��  �<  #0w0  2�:  ?1�  2	�  ?
  �  �  G  T3%  "4�'  3�5I  s   �  �  6�  7{�  �  	:�  8tR    9��  P%   M 3
  !� :�  #;Z�  �%  ��  ��  !�  #�S   �  %3_  %�  '<j�  �  x  ��  ��    %�  &��  '=՘  (�l  *�  +2�  $�A  +�� �ڇ   UW    �  #�  $	  %'	  7	  &P	  `	  '>7  4  (�	  �	  �)�  *M6  �#  +��  ,P'  -`'  p'  	.��  �'  y/��  !iN    �<  #0w0  2�:  ?1�  2	�  ?
  �  �  G  T3%  "4�'  3�5I  s   �  �  6�  0  �z  	{�  
W�  x�  7��  ?8��  9�  �  �r  �  :�  :tR  ;��  P%  "��  ��  ��    �%  $3_  �  &  !�S  f   <Z�  "��  ��  %�  '=j�  �  x  "%�  &��  '>՘  (�l  *�  +2�  ! �A  -�� 4�   �`    �  !�  "	  #'	  7	  $P	  `	  %>7  4  &�	  �	  �'�  (M6  �#  )��  *P'  +`'  p'  	,��  �'  y-��  iN    �<  #.w0  2�:  ?/�  0	�  ?
  �  �  G  T1%  "2�'  1�3I  s   �  �  4�  	x�  5��  ?6��  7�  {�  �  �r  
�  :�  8tR  9��  P%  "��  ��  ��    �%  $3_  �  &  !�S  f   :Z�   ��  ��  %�  'j�  �  x   %�  &��  ';՘  (�l  *�  +2�  !�A  ��� �a�   �o      ��  ��  x�  �  �  	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  ��  ? ��  �<  #!w0  2�:  ?"�  #	�  ?
  �  �  G  T$%  "%�'  $�&I  s   �  �  '�  ({�  �  !	�  #�S  
�%   �  %3_  %�  ')j�  �  x  ��  ��    &  (*tR  +��  P%   �A    �s    �  %�  &	  ''	  7	  (P	  `	  )>7  4  *�	  �	  �+�  ,M6  �#  -��  .P'  /`'  p'  	0��  �'  y1��  ˈ  �<  #$w0  2�:  ?2�  3	�  ?
  �  �  G  T4%  "5�'  4�6I  s   �  �  7�  8�  9��     	x�  :��  ?;��  <�  {�  �  =�9  #iN  
  >�  0   �z  W�  "?Z�  #�  '  2  @��  ��  !�  #�S   �  %3_  %�  'j�  �  x  ��  ��    (A3  @%�  &��  '"՘  (�l  *�  +2�  $!�r   :�  f  (\� )"�   #�     �  �  		  
'	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  !��  P'  `'  p'  	��  �'  y��  "��  ?��  #;�  %�9  &��  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  T�� U�� V�� W�� X� Yώ Z�� [� ]� _8� c'� ��� �X    �� �� ��   �    ��  P'  	  '	  7	  	P	  `	  
`'  p'  	��  �'  y��  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  K � � o�� q%�   Y�    �  �  	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  ��  P'  `'  p'  	��  �'  y��  ��  ?��  ��  ��  x�  �<  #w0  2�:  ?�   	�  ?
  �  �  G  T!%  ""�'  !�#I  s   �  �  $�  %{�  �  &��  	  
�%  $3_  �  &  !'�S   (�  &)  (*tR  +��  P%  @  ,�
 8�   q�    �  $�  %	  &'	  7	  'P	  `	  (>7  4  )�	  �	  �*�  +M6  �#  ,�  ˈ  �<  #-w0  2�:  ?.�  /	�  ?
  �  �  G  T0%  "1�'  0�2I  s   �  �  3�  4�  5��     x�  6��  ?7��  8�  9{�  �  	0  �H  
j�  "�  :�9  #iN    ;�   �z  W�  "&�  �    #w� ��    !�  #�S  �%   �  %3_  %�  �  $<Z�  =��  x  ��  ��    (>3  =%�  &��  '?՘  ( �l  *!�  +"2�    ��    �  2�  3	  4'	  7	  5P	  `	  6>7  4  7�	  �	  �8�  9M6  �#  :iN    �<  #;w0  2�:  ?<�  =	�  ?
  �  �  G  T>%  "?�'  >�@I  s   �  �  �  	�  
0  0X{  7  / �z  {�  W�   ˈ  A�  B�  C��     !D�@  "x�  E��  ?F��  G�  �  #H@  %| '&�  �    (w� ��    !�  #�S  �%   �  %3_  'j�  �  )IZ�  J��  x  ��  ��    (K3  J% �  &!��  'L՘  ("�l  *#�  +$2�  +%�  �&�  ,1�l .'#  1*� )K (� 4+V  7-�r  ,:�  f  :.#�  Mw  #  D�� E�� F#� G� I�� M@� P@� S�� T�� VJ� W͗ [� ^,� _�� `ĕ a<� c>� f� h�� k� lT� m�� nߓ o� p'� rl� s�� u�� vT� w(� x#� y˚ {ߖ �� ��� ��� ��� ��� ��� ��� �Ù �� �� �� �!� �i� ��� �O� �� ��� �� �֕ �� �� �� ��� ��� ��� ��� �n� �z� �ޙ �|� �^� �A� �{� �+� �Й �^� �і ��� �ǝ �Y� �'� �'� �x� �h� �� �G� �y� ��� �� �Л �ܜ ��� �� �;� ��� �� ��� �"� �l� �9� �� �� �X� ��� ��� ��� ��� �� �I� �=� �� �:� �Ô ��� �Ҕ ��� �� �z� �^� ��� ��   ��    �  (�  )	  *'	  7	  +P	  `	  ,>7  4  -�	  �	  �.�  /M6  �#  0��  1P'  2`'  p'  	3��  �'  y4��  � �<  #5w0  2�:  ?6�  7	�  ?
  �  �  G  T8%  "9�'  8�:I  s   �  �  &iN    ;�  <�  =�  �r  ��  
x�  >��  ??��  @�  	{�  �  %  :�  AtR  B��  P%  "��  ��  ��    �%  $3_  �  &  !�S  f  K � !'X{  -  "C #@  %!��  DZ�  E��  ��  %�  'Fj�  �  x  E%�  &��  'G՘  (�l  *�  + 2�  �  �"�  &$�z  #W�  '%0  ,p� 4�� 8�� <ğ >)� ?�� @�   5�    !#�  %�<  #w0  P	  	`	  2�:  ?
�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  '  2    2�    �  �  	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  ��  ?��  �?  iN    �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  " �'  �!I  s   �  �  "�  #Ə  $�  A,  %�9   �  !M &  "X{    #	�H  j�  "�  $�z  '{�  
W�  %0  '(w+  .��  �ܡ �;�   j�    �  +�  ,	  -'	  7	  .P	  `	  />7  4  0�	  �	  �1�  2M6  �#  0  )X{  0  �<  #3w0  2�:  ?4�  5	�  ?
  �  �  G  T6%  "7�'  6�8I  s   �  �  * ˈ  9�  :�  ;��     <�9  =iN  	  
�  �z  {�  W�  !| x�  >��  ??��  @�  �  #AZ�  #�  '  2  B��  ��  !�  #�S   �  %3_  %�  'j�  �  x  ��  ��    (C3  B%�  &��  'D՘  (�l  * �  +!2�  $$� #K "� &&�r  %:�  f  ,'V  .(� =�� >�� KQ� L�� O� P� R�� S� W�� X5� Z�� ^ � _g� a� c�� e�� fa� gʥ hU� �r� �� �s� �� ��� ��� ��� �� ���   ��    �  �  	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  
��  P'  `'  p'  	��  �'  y��  ��  ?��  X{    �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  ��   $ 	�z  !{�  W�    
�    �  	�  
	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  w+  �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  @  W�    %�    �  
5�  {�  �<  #w0  P	  `	  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  c,  @  c ��  	�z  �  �  	  '	  7	  >7  4  �	  �	  ��  M6  �#  W�  0     K� V� 5�   ��    �  �  �  	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  ��  P'  `'  p'  	��  �'  y��  ��  ?��  �<  #w0  2�:  ? �  !	�  ?
  �  �  G  T"%  "#�'  "�$I  s   �  �  %w+  5�  {�  c,  &�9   iN  '  (�  !�  "X{    #	0  %�z  
W�    }�    	�w  �  
�  	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  E�s  iN    �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  �  $�� %� ��   �     �  
�  	  '	  7	  P	  `	  >7  4  �	  �	  ��  M6  �#  	X{    �<  #w0  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  W�  0        ��  P'  	  '	  7	  P	  `	  `'  p'  	��  �'  y��  �  �?  ��  ?��  �� ��   �  !�  "�] 	#M6  
$*F f�  �  %>7  4  &�	  �	  �'$�  (w+  )Ə  *�  A,  �<  #+w0  2�:  ?,�  -	�  ?
  �  �  G  T.%  "/�'  .�0I  s   �  �  1@  2�2  3iN  4  �  5�9  6�   �  !	�� "
@  #��  $7X{  &  %#�  '  2  &�H  8j�  "�  '�z  9{�  W�  (:0  *�V     �� &� � � �� 	i� 
� ,� �� 
� �� � ?� Ь ٫ {� � �� ��    ~� �� �� �� �� 	K� 
Ƭ V� ϫ |� �� %� �� �� �� ��    Y� � ܰ � +� 1� <� �� �� �� � `� ϭ h�  �� !Y� "� #�� $ʯ (U� )� *D� +ͮ ,� -� @�� AE� Bq� C�� DY� F�    �  �#    �	    w+  �H  �<  #w0  P	  `	  2�:  ?�  	�  ?
  �  �  G  T%  "�'  �I  s   �  �  j�  "�  @  �   
� 	x�  �  �  	  '	  7	  >7  4   �	  �	  �!�  "M6  �#  #��  ?$��  %�  &{�  �  !�  "0  $#�  '  2  %'@  '�V  )(�  *��  )P'  *`'  p'  	+��  �'  y,��  ,-�� .��  /�  0�] 
1*F f�  .   02B^ 	3�` 
4�J 5�D 6�a 7�a 8Na 9�] :�] ;�] <Q` =.^ >P^ �� �k� �̲ ���    �� !O� "2� #� 4��   �    eK 	�  ?
  �  �  u�     5K  K   � i�   �  �  	  '	  =�  P	  `	  >7  4  �	  �	  ��  M6  �#  V�  l�  	�  ��  �  �  *3  	�  
s� 	 �� ��  ?!��  �  "� $
)!�  �"��  �##� ��  Q�  K��  $P'  %`'  a�  	&��  �'  y'��  La� M��  ��  (��  6�  �  	Ѹ 
>� � � d� C� )@  �V      .%   q�  #'   
   �5       h   �&   =   �
   �   3*      +7   �%   �:   �   �!   �    �   ,   �%   ?2   ?   Z$   w&   �   �   x5   >>   m      K,   >	   �(   O3   T�  e   �<   B   �%   �   	+   o   �   MB   �0   n   �   �7   V2   �    e1   R   �   �      �	   �   �   �   �9   �'   �<   J&   �   �0   �4   	   ?A      $   �5      ��  8�  ��   �  ��  ��  o�  ��  �  ��  B�  `�  (�  |�  ��  ��  ��  ��  $�  �  ��  ^�  m�  ��  ��  ��  `�  3�  �  ��  x�  �  �  '�  .�  P�  u�  ��  S   T
   �+   �   �.   �   4   �	   1   �&   �   t:   #&   s2   O4   z6   �   �   6-   �@   �5   0�  ��  �   0   �8   I/   ;   ;    1(   �+   U   �%   	*   v*   ^   q       �6   �   �   G   "
   /$   1   
A   �0   �8      �;   +   �   �&   �   F*   �?   5&   )#   F   �-   	C   ;   Y   t   �2   B   �C   �   �)   �!   �   4    0   �   2   (   �   t;   �   �   04   K   ?   (   7   �   �,   �   �7   :;   1   C   �$   p   \   �   *      k%   �=   �    u�  ��  ��  |�  �	   �;   �   '   �   -   j   �   pA   �C   `4   �    e	   5'      �      �0   w   �   L   �	      �@   �   �   �A   .   Z)   =
   �   ^   SC   �
   t<   �      T      P"   �   d3   r@   �   k   Y    �   �   B   �(   �   O   �@   �   j   �1   W>   �B   x   �.   �    Q    0   /   �   �?      �   �#         �   ^   �=   �3   �         �   !   �:   e   c-   J   eB      �/   �$   5)   z7   0   �   O   �   m$   iC   �   �.   �A   -   �   `/   �      :+   �/   Z?   H-   �<   �?   �%   �=   �   )   g      �!   �=   y   ;5   ,   �:   ~   3    �6   �   x4   >$   1B   �   �(   �   �   @   H   V.   �   �=   5   �5   �   #   �6   !   �   �   >   9%   �8   �*   �2   �4   �*   �9   �   �#   -;   �!   �     ��Q  �ݶ ��     �� >� �    � �� �� D�    3  �  �  �   W  "�  #�,  $�  %  (�  )�&  *�/  +>  -E  .:  /�  0S  2�  3�+  4$=  5P@  R�>  S  T�+  W<  X*  Y�  \    ]R+  ^  a�  b$6  c^(  �I:  ��  ��;  ��  �O7  ��3  ��  �$  ��9  �.  ��,  ��4  �  �t
  ��  ��>  �\8  �x  �F=  ��  ��#  �W0  ��1  ��  �>8  ��  �c   �G� �3     �� *� h� � 	� 
l� �� � L� �� �� �� �� � �� 8� O� }� �� �� e� �� �� �� ,� � $�  �� !�� "�� #�� $7� %{� &�� '�� (�� )� *ý +9� ,�� -�� /��    '�� (�� *�� �[� �T� �)� �j� �>� �:� �Q� �W� ��� �� ��)  ���  ���  ���  ���  � �  �.�  ��  ��  ���  �W�  ���  �u�  ���  ���  ���  ���  ��  ��Q  �ݶ ��  �4� ��� �a�    �� "�� %� .�� 2S� 6˼ C�� F�� R�� V�� ^X� c�� l�� m� vӽ �k� ��� ��� ��� ��� �(� �b� �� ��� ��� ��� ��� ��� ��� �q� ��� ��� ��� ��� ��� ��� ��� ��� �s� �� �x� �s� � � ��� �r� ��� �� ��� ��� �Y� ��� �S� �־ ���    �� '�    �^� �(� ��� �+� �K� �� ��� �min �max ��� �� �� ��� �� �N� ��� �1� �� �j� �� ��� �� �Q� �M� �5� �� �s� �÷ ��� �w� �b� �Ŷ �"� �r� ��� �� �,� �%� ��� �S� �7� �~� �K� �{� ��� �>� �_� �� �� �� �n� ��� ��� �~� ��� ��� �3� �U� ��� ��� ��� ��� ��� ��� ��� �ٷ �s� �� �X� ��� �&� �t� ��� ��� �b� �h� ��� �� �K� �Ͽ �'� �e� �� �0� �� ��� �� �� �� �>� �� �	� �8� ��� ��� �
� ��� �� ��� �N� ��� ��� ��� ��� �4� ��� �$� ��� ��� �x� ��� �� ��� �� ��� �K� ��� ��� ��� �=� �� ��� �`� ��� ��� ��� ��� �ڻ �E� ��� ��� ��� �� �
�� �
5� �
� �
�� �
�� �
�� �
�� �
��  �
�� �
�� �
�� �
�� �
f� ��� �L� ��� �h� ��� �M� �� �d� �{� �W� �g� ��� ��� �c� ��� �z� �� �� ��� �� �:� ��� �� �>� �w�    ,~� J��    �� ��)  ��  ��Q  �ݶ ��  �4�    /� %�� *a� ,abs    P��  T�� WZ� Z�M [� \�� ]�� ^� _div `c� am�  b� c2� d� e��  f�� gN� h�� i�� l]� o� p�� q� r�� s� t�� uC vl� w�� ��� �1� �� ��� � � �_� ��� ��    �� P� � e� � |� F� 	� 
N� h� M� f� �� '� Ѹ >� � � W� g� H� � �� �� ��    �� 8� G� � 	�� 
�� 7� 9� W� ,� �� ��                                      X@                   h@                   �@                   �@                   (@                   X@                   0@                   @@                  	 �@                  
 �JB                   �JB                   ��C                   0Yd                   8Yd                   HYd                   XYd                   �Zd                   �Zd                   @\d                   ��e                                                                                                                                                                                                                                                                   ��                     8Yd                  HYd             (     �C             ;    	 0@             =    	 `@             P    	 �@             f      �e            u     �e            �    	 0@             �      �e     0           ��                �     @Yd             �     (YD             �    	 `JB             �    ��                �    ��                �    	 /B     �       �     -f                 -f             #    -f            <   	 @            R   ��                Z   ��                �    ��e            c    ��e            g    x�e            �    ȕe            �    ��e            �    ĕe            r    ��e            v    ��e            {    ��e            �    ��e            �    ��e            �    ��e            �    ��e            �    �\d            �    p�e            �    �\d            �    ��e            �    ��e     P       �    ��e            �    ��e            �    ��e            �    ��e            �    ��e            �    ��e            �    ��e                ؕe                ��e            B3    �e                ��e                �e            (    ̕e            5    Еe            B    p\d            Q     �e     P       Z    ��e            ^     �e            b    P\d            t    �\d            q    D\d            �    @\d            �    ��e            �7    �e            �    ��e            �    �e            �    ��e            �    ��e            �    `KB             �    ��e            �    ��e            �    p�e            �    @KB               ��                    $�e            #    @�e            *     �e            4   ��                =   	 �&@     K       G   	 
'@     #       X    @�e            \    `�e            f    �PB     P      l   ��                u   	 �*@     ?       �    ��e             �   	 �*@     .       �    X`d            �   	 �*@     �       	    ��e            �    Пe            �    ��e      P      �    ȟe            �    ̟e            �    ��e            �    d�e            �    ��e                h�e                p�e               ��                !   	 .0@     K       *    \`d            <    ��e            Q    ��e            a    ��e            y    ��e            �    ��e            �    �\B     0       �    �\B     �       �   ��                �    �^B     �       �    `^B     P       �     ^B     H       �   ��                �   	 �D@     �       �     �e     P           �`d                ��                #    �ad     �      /    P�e            >   ��                G    `�e            P    h�e            �0    X�e            ]    p�e            l    x�e            o    �B     0       z   ��                �     �e            �    ��e     $       �    @�e     T       �    ��e            �    ��e            �    ��e            �    ��e            �    ��e            �     �e            �     �B     H       �    ��B     @       �    ��e                ��e                ��e            #    ��e            /    ��e            8     �e            E    ��e            P     �e             `    ��B            k    ��B     0       v    ��e            �    ��e     P       �   ��                �   ��                �     �e            �    �e            �    @�e     �      �    �e            �    p�e            �     �e     p       �    `�e     �       �     �e                D�e                $�e                 @�e            �E    ��e            1e    |�e            *    ��e     �       4    x�e            A    t�e            U     �e     Q       f   ��                q   ��                ~    ��e            �    �7e     (       �    �7e            �    ��e            �    �7e            �    �7e            �    ��e            �    |�e                x�e            #   ��                -    ��e            :    ��e            G   ��                R    ��e            ]    ��e            n    �7e            }    h�B     
       �     8e            �    X�B     
       �    H�B     
       �    ��e     
       �   ��                �    ��e            �   ��                �   ��                �   ��                �   ��                	   	 8�@     F       	   	 ~�@     F       &	     Ge            4	     8e            C	   	 ď@     9       U	    ��e            i	    ��e            ~	    ��B            �	    @8e     �      �	    @Ge     �	      �	   ��                �	   ��                �	   ��                �	    �B            �	    ЧB            �	    ��e            �	    ��e            �	     �e            �	    ��e            
    ��e            
    ��e            %
    ��e            0
    ��e            <
   ��                E
   ��                P
    �B            Y
   ��                d
   ��                n
   ��                x
    �e            �
   ��                �
   ��                �
   ��                �
   ��                �
    �e            �
   ��                �
   	 5A     t       �
    @�B     (      �
   	 �A     1          ��                     �e     �          ��                )   ��                2   	 �.A            ?   ��                I   	 t:A     R       V   	 �:A            d   	 �:A     -       r   	 ;A            �   	 ;A     ^       �   	 };A     +       �   	 �;A     Q       �   	 �;A            �   	 <A     7       �   	 H<A     )       �   	 q<A     &       �    �e                �e                 �e            '   ��                1    ��e            Q     �e     �       b    ��e            m   ��                w   ��                �    �[e            �    ��e            �    ��e            �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �    ��e               ��                   ��                   ��                (   ��                0   ��                ;    ��e     �      C    @f     �      K   ��                R   	 ��A     +      \   ��                g    �f            k    �f            z   ��                �   ��                �   	 0�A            �   	 C�A     `      �    �$f     P       �    �$f     P       �    �$f            �    @$f     0       D    �"f            5    `"f     `       M    �"f     P      �    �"f            �    0%f            �   	 ��A            �    H%f                 X%f                `%f                 f     4           �e            *    �f            8    �f            F    Lf            S    Pf            `    `f     $       p    h�e            }    �e            �    8f            �     �e            �     "f     0       U    @f            �    �f            �    @%f            �    <%f            �    8%f            �    L%f            �    P%f                4f                T%f                `f     �            �f     �       *    �!f     8       3    @ f            :     f     8       B    `!f     0       K      f     0       S    `f     �       ^    �!f     0       f    D%f            q    �e            |   ��                �   	 ��A     8       &$    x%f            �   	 &�A           �    t%f            �    h%f            �    p%f            �   ��                �   ��                �    �%f            �    �%f            �   ��                
   	 hB               	 {B     @      ,    �'f            5    0&f            <    �&f            D    �'f            H    p'f            L    `'f            R    @�C            [     �C             a    @�e     �      �     'f     P       �    X'f            o    �&f            x    �&f            ^    �&f            �    �&f            �    �&f            T    �&f                �&f            �    P'f            �    �&f            �    �&f            y    �&f            �    �&f            �    �&f            �    �&f            �>    `&f             �    @&f             �    (&f            �   	 �B            �    `�C            �    �'f            5    �'f            �    �'f            �    �'f            �    $&f                �'f                 &f                �'f                �%f     @       "    �%f            �>    �'f            ,    �&f            -    �&f            2    �%f            ;    �%f            E    �'f            P    �'f            Z    �'f            d    �%f            l    �%f            u    �'f            }    �'f            �    ��e     �      �    ��e     �      �   ��                �    �'f            �     (f            �   ��                �   ��                �   ��                �    (f            �    `�C     @       �   ��                �   ��                   	 Q)B               	 g)B     P       )   ��                3    (f            =    ��C     �       H   ��                R    @(f            Y    @,f     4       ^   ��                l   ��                t   ��                �   ��                �   ��                �    	 �HB             �    	 IB             �    	 MIB             �    	 WIB             �    	 �IB                 	 �IB                ��                "   ��                -   ��                4   ��                =   ��                G   ��                Q   ��                Y   ��                d   ��                     ��                n    XYd             w    �Zd             �   	 (�@     W      �  " 	 �EB     -       �    P-f            �    �6f            �     (f            �   	 �@     -       �   	 i
B            �    `Df            �   	 \bA     �          	 f�@     >          	 ~A     "         	 �1B     8       6    @zg            E    �ef            P    @Xe     (       W   	 "�@     p       l   	 1�@     5       �    �6f            �    @Re            �    �Pe            �   	 �@     K       �    (ce            �   	 H�A     �       �   	 r+A     �      �   	 �%@     t       �    �Pe            �   	 ��A     �       �    ��e            �   	 ~eA     6           `-f            
    ��i               	 	�@     :       *   	 ��@            5    `If            E   	 ݛA     �       \    �6f            d    T�e            y    hDf               	 ��@     -       �   	 �CB     �       �   	 )�A           Y    �e            �   	 �&B     �       �   	 ѹ@            �   	 {�A            �   	 hA     |            �i                �Pe               	 ��A     �           lDf            #                     *   	 �@            I$    `_f            7    p6f            @   	 �<A     8       S   	 2�@     �       `    pDf            f    ��i            t   	 �/A     M       �   	 ob@     V       �   	 =�A            �   	 �@     +      �   	 �~@     �      �   	 �@     .       �  " 	 �GB     -      �   	 ��@            �    p[e               	 ��A     �           ��B      �          	 �~@            (   	 -9A            1   	 OA     
      G   	 J�A            X   	 A     �      d     Ve             n                     v   	 :�A     /       �   	 `�A            �   	 C9A            �    ��f            �    ��f            �    |Qe            �   	 ��@            �    ��f            �   	 89A            �   	  A     �       �    تf            �   	 �B           	   	 	2@     R           Bf            *    �Qe            6   	 \IB             D    �Qe            P    tDf            b    �Qe            n    �7f            v    �_d     �       �   	 ��@            �   	 ��@            �    �7f            �   	 8@     J       �   	 ��A           �    xDf            �   	 4B     �      �   	 Ɵ@     "       �    �`f               	 �S@              " 	 �EB     -       -    hIf            6    �Qe            A   	 o"B            Q   	 )*@     0       c   	 �@     T       v     Hf            �     Re            �   	 �s@     X      �   	 �.B            �   	 D�@     H       �   	 JeA     4       �   	 4A     �       �    pIf            �    |Df               	 /0A     _         	 ��@     �           ��i            )   	 ��@     6       C   	 �B     6       R   	 zHA     �      f   	 �W@     	       t                     {   	 8�@     i       �    �e            �   	 ��@            �   	 �WA     �       �    ,Qe            �   	 2�A            �    �~e     �      �   	 �A     z       �   	 [~@     3       �   	 � A           	     8f               	 �U@     �           	 �0B            +    �Df            6   	 ,A     �       E    `}g            N    T-f            W   	 �@     p       f     Qe            w   	 �A     e       �   	 v�@     #       �    $Qe            �     �i            �   	 �@     g       �   	 ��@            �     9f            �   	 �A     ]       �    �We     �       �   	 	�@     R          	 � @     �           9f            *    ��f            6    �ed            B   	 *�A     �       M   	 �C@     '       ]   	 -B     /       f   	 �/@     /       z    �Df            �    �Re             �    �Qe            �   	 qj@     7      �   	 A�@     5       �    d-f            �    9f            �   	 k�@     I       �   	 �A     b       �    x6f            �*                     �   	 ��A     �          
 �JB                	 �@     $          	 �9A     $       -   	 {"@     s       7    ��C      @      C   	 �>B     >       XF     ed     �       b   	 4B     .       l     Df            s  " 	 �DB     �       �   	 !U@     �       �    �Jf            �    �i            �   	 ��@     �       �   	 x8A     �       �    �Df     P       �   	 �#B     7       �    �`f            �  " 	 �DB     2          	 �k@     �         	 TxA     �            Ye     (            �f            5   	 A�@     �       <    9f            H    �Pe            X   	 f*B            d  " 	 vEB            s    TRe            |   	 <q@            �    ��g            �  " 	 JB            �    �Qe            �    tQe            �   	 �A     �      �    �6f            �   	 �A            �                     �    xQe            �   	 �.B               	 ١@     4       %   	 �A            <   	 �_@     �      H    ��i      (      S   	 E+A     -       c    0Qe            q    pQe            }   	 ��A     A       �    9f            �   	 �A     m       �    ��f            �    �Re     �       �   	 ��@            �   	 �@     6       �    �`f            �   	 �c@            �    ��i     �      �    �`f            �   	 ��@     �           �f                 h_f            (    	 /.B            5    	 �&@     2       @    	 O3B     u       f    	 �@     /       r    	 �1@                	 �A     s       �    	 �TA     �       �     ��i            �    	 O�@     �       �    	 �}@            �    	 ~�A     �       �     9f            �    	 ��A     N       �    	 W�A           !    �Qe             !   	 
�@     A       *!   	 �kA     $      5!    �Se     �       >!   	 3A     >       F!    �gf            R!    tIf            [!    0Df            e!    9f            u!   	 4&B     P       �!   	 ~B     |       �!    �_f     d       �!   	 �aA     �       �!  " 	 �IB     )       �!   	 ��A            �!    �ed            �!   	 � B            �!   	 IB             �!   	 .vA            �!   	 �^A     s       "    �f            "   	 �vA     x       #"    ��g            /"    ��f            7"    (Hf            A"   	 m�@     9       O"    ��e            X"   	 �i@     `       d"   	 ߚ@     #       r"   	 A�A     �       z"   	 I8B     j      �"   	 W5A     &       �"   	 �#@     �       �"   	 &�@     R      �"    ��f            �"   	 ��@            �"   	 �O@            �"   	 ��@            #    @�i     �      #   	 sQ@     _      )#   	 �A     
       9#    xIf            =#   	 >A     �       I#    ��f            V#    �i            _#   	 t}@     4       o#   	 ��A     �       #    ��e            �#   	 �A           �#                     �#    ��g            �#   	 ��@            �#    |If            �#   	 �/B     E       �#    ��f            �#    ��f            �#    �`f            �#    �Jf            �#   	 �o@     U      $   	 A�@     b       $    �\d     H       "$    l�e            /$   	 �+@     `       9$   	 �5A     R       F$    �_f                 �_f            T$    �If            X$    �Ze             _$   	 �B            �E    �_f            q$    ��f            w$    ��f            �$   	 �y@            �$   	 ڿ@     u      �$    Bf            �$    ��e            �$    ��f            �$   	 ^B            �$   	 [&@     2       �$   	 �`A     �       �$   	 �1A            �$   	 &%B           �$    ``d            %   	 1B     1       +%                     2%   	 h�A            A%    �Qe            X%    �Df            a%                     i%   	 �9A            t%   	 z@     *       �%    ��g            �%                     �%    �jd     P       �%   	 ̙@     :       �%    ��f            �%    (Df            �%    `be     �       �%   	 �P@     �       �%    PRe            �%    9f            �%   	 �@B     C       	&   	 �A     q      &    @_d     @       '&   	 {@     �       ;&   	 v�@     �       M&    �Pe            w2    �If     �       \&    ((f            m&   	 M4B     I       �&   	 &�@     e       �&                     �&    �i            �&    �`f            �&   	 ݆@            �&     ]d     0       KZ    ��f            �&   	 �A     }       �&   	 4(A     [       '   	 N9A     �       '    �i            "'   	 �qA     �      fS     9f            3'    ̓e            C'    �i            R'    HRe            a'    `�e            l'   	 �@     �      {'   	 �,@     :       �'    �Qe            �'                     �'    ��f            �'   	 �6A     m       �'    <Qe            �'    ��i            �'    (9f            �'     �g            �'   	 {pA     Z      (   	 ��@     !       (   	 ��@     �       (    d`d            ((   	 dH@            6(   	 ��A           E(   	 Az@     #       _(    �e            m(    x�e            x(   	 �@     B       �(    ��e     H       �(    �i            �(   	 I�@           �(   	 ��@     �       �(   	 +6@     �      �(    ��B            �(   	 �}@     #       �(  " 	 �EB            )   	 �3B     [       #)   	 B�@            .)   	 �@     >       ;)   	 _�@     �       H)    ,9f            Q)   	 �eA     F      [     af     �      d)   	 ��@            s)    �Df            z)   	 -�@           �1    ��f     �      �)   	 eA     5       �)   	 (?A     �      �)   	 �@             �)    0Hf            �)   	 ��@     )       �)    h-f            �)   	 �@     1      �)   	 �0B     2       �)   	 k�A             
*   	 �A            *                     !*   	 �2A     /       **    @_f            5*   	 �0B     $       G*   	 �"B     K       X*   	 w�A     e       f*   	 ȳ@     >       s*   	 +�@     R       �*   	 ��A     �       �*     �i            �*     Re            �*   	 �-A     .      +    09f            �*   	 �@     �       �*    �Ze            �*   	 [�@            �*   	 �0@     .      �*   	 X-B            	+   	 dI@           +    49f            "+   	 �9B     W       X+    Re            a+   	 ��@     S       p+   	 �$@     d       ~+    89f            -_   	 �@     	      �O    0@             �+    ��e            �+    �ed            �+   	 iA     W       �+   	 �cA            �+   	 �@     �       �+                     �+   	 ˂@     %       �+   	 3A     b      ,   	 ��@     D      ,    �ed            #,    ��f            /,   	 B     �       >,   	 ��@     �       N,    @9f            U,   	 ]@            j,    ��f            u,   	 _A     �      �,     �f            �,   	 �"A     2      �,    �Df            �,     �g            �,   	 5A     �      �,                     �,   	 �D@            �,   	 �.B            -   	 ~�@     +       -   	 w�A     �       *-   PYd             7-    4Re            A-   	 ��@     9       S-    @Jf            [-   	 lB     
       i-   	 �@     ]       r-   	 ��@     +       |-    �Ue     (       �-   	 ��A             �-   	 �A     e      �-   	 �1A            �-    8Re            �-    �Df            �-   	 ��@            �-   	 �(B     ,       �-   	 އ@            �-    `Ue     (       �-   	 vA            �-    HJf            �-    t�e            .   	 �%@     %       .   	 �@     J       &.   	 ��@     �       -.    $(f            >.    ��e     H       M.   	 �B     n       W.   	 Z6A     e       a.    �_f            n.    $�i            v.   	 {	B     /       �.   	 
}A           �.   	 ��@     4       �.    8Hf            �.   	 F'B     �       �.                     �.    Re            �.    �Jf            �.   	 9^A     h       �.   	 B            �.   	 �"@     �       /   	 ��A           /   	 �4B           5/    �7e            C/   	 ��@     6       T/    4Qe            b/    �^d            n/   	 �W@     Q      |/   	 ��@     
       �/    PJf            �/    H9f            �/                     �/  " 	 �FB     "       �/    �Pe            �/    (�i            �/   	 �v@     ;      �/    hQe            �/  " 	 �DB     2       0    `Qe            0   	 �<A     �       0   	 i�A     �      *0    ��f            40    �Df            ?0   	 dA     7       ]0   	 ��A     ,       l0     Wf            u0   	 �	B     �       �0   	 �@     E       �0   	 X@     1       �0    �`f            �0                     �0    @�f            �0    Pif            �0   	 �.A     �       �0   	 �A     L       �0   	 �AA     �      �0   	 ��A            1    �Jf            1   	 +|@     Z       #1   	 '$B     T       *1   	 4�@            =1   	 �.B     I       O1    TJf            Z1   	 un@     �       f1   	 �A            u1    LQe            �1    P9f            �1   	 b�A            �1   	 �@     Y       �1     �f            �1    �`f            �1   	 #�A            �1     Ef            �1   	 ��@     �       �1    �f            �1    �Pe            �1     `f     (       2    l-f            2   	 YA     �       (2   	 Q?B     /       =2    (`f            J2    �ed            T2    XJf            _2    �6f            g2   	 ��@     &      t2    `Jf            2    �Qe            �2   	 k�@     B       �2   	 Oj@     "       �2    �Qe            �2    �Ze            �2   	 0�@     +       �2    p-f            �2   	 ��@            �2   	 vB            �2   	 8D@     -       �2   	 �@     �       3   	 YA     ?      3    �7e            +3     Gf     �       :3   	 �*B     �       E3   	 NA     z       T3   	 ��A            d3   	 �@     �       u3    Re            �3   	 �FA     �      �3   	 }@     U       �3    �f            �3   	 g*B     a       �3   	 ��A     �       �3   	 ��@            �3    x-f            �3   	 7�@     .      �3   	 �tA     �      4    0�i            4   	 ܛA            &4    �7e            34    (f            <4    dQe            I4    �Ue             S4   	 �{A     �       j4    X9f            u4   	 �|A     Y       �4    PQe            �4   	 ��@     e      �4                     �4   	 ��A     A      �4                     �4   	 �A            �4   	 �.B            �4    0`f            �4   	 DdA     �       �4   	 �O@     �       5   	 PB     W       5   	 9�@     �       -5    @ce     @      35    �-f            <5   	 �5A     e       J5   	 �A     m       \5   	 >.B     ]       i5    pJf            p5   	 ��A     !       5   	 r�@            �5   	 JS@     ^       �5   	 �mA     �      �5   	 �'@     �      �5   	 p�@            �5   	 Y*@     5       �5   	 ��@     �      �5    \9f            �5    �-f            �5   	 eiA     �       6   	 Y-B     �       6    Re            +6    �Qe            96     �i            �   	 ��@     �      K6    �Qe            X6    �f            c6    �Qe            t6    D�f            �6    �Jf            �6    �Qe            �6   	 H�@            �6   	  6@            �6   	 ��@            �6    �7e            �6   	 ��@     $       �6   	  �@            �6    `�e     H       �6   	 ��A     :       7    �Qe            7   	 (�@            7   	 ��A     �       07   	 ,�@     D       A7    �Re     (       I7   	 ��A     )       R7   	 �;B     �       v7   	 �SA     �       �7   	 �AB     �       �7   	 �)A           �7   	 `�@     �       �7    �f            �7   	 �#A     L      �7    `if            �7    ��i            �7                     �7    HQe            8    �Qe            8   	 7%A     �      !8    8�i            .8    �6f            :8    `9f            g    8`f            �    �-f     �       F8    H�f            T8    d9f            [8   	 s�@            l8    �Jf            u8  " 	 �FB     �       �8   	 �7@     �      �8   	 ��A     q       �8   	 j�@     h       �8   	 �f@            �8    h9f            �8    Ef            �/                     �8   	 ��A     q       �8   	 �1B     �       9   	 �@     "       !9   	 �A     �       /9   	 b@     #       D9   	 �.B            U9    @`f            ^9   	 i(B     V       k9   	 �B     2       v9    Qe            �9    �if            �9   	 B            Y    �f            �9    �`d            �9   	 5�A     G       �9   	 ː@            �9   	 �@     R       �9    @-f            �9     �g            �9    @�g            �9                      :   	 �A     �      :   	 F�A     �       !:   	 �A     �       6:    x,f            F:     Ve     (       Q:   	 �@     B       e:    XQe            u:   	 �A            �:   	 ~@     ?       �:   	 �A     #       �:   	 )�@           �:   	 �.B            �:    L�f            �:    p9f            �:    �Qe            e   	 @            �:   	 ��A     1       �:   	 g@     }      �:    �Jf            ;    ȴi            ;    �Qe            !;    <�i            (;    P�f            2;   	 �(A           A;    @�i            K;    <Re            S;    X�f            ^;   	 ��@     �       i;   	 �B     �       ;    �f            �;   	 D�A            �;    D�i            �;   	 BcA     .       �;     Qe            �;   	 }�@            �;   	 �A     �       �;   	 �@     �       �;   	 ��A            �;    `�f            �;    �f             <    `�f            <   	 e�@     �       !<   	 VvA     E       /<    дi            <<   	 �B     v       M<    t9f            [<   	 �~@     F       c<                     k<   	 ��@     Z       x<    �if            <   	 wA     B       �<    �Jf            �<    �Jf            �<   	 d�@            �<    Ef            �<    �6f            �<    $Re            �<    DQe            �<   	 pMA     �      �<   	 �"B            =    D`f            =   	 UwA     �       =   	 dz@     �       0=   	 �!B     �       ?=   	 L�@     *       Q=    H`f            Z=   	 �@     :       i=    d�f            q=    �hd     h      z=    شi            �=                     �=   	 �|@     D       �=    �Qe            �=   	 �|@     V       �=   	 Is@     ;       �=    �f            �=   	 5�A     &       �=    �Qe            �=    �i     ,      �=   	 8SA     �       	>   	 �A     +      >    �%f            >   	 O�A           0>    �Qe            =>   	 x�@     #       L>   	 EA     	      ]>    Ef            g>   	 ��@     x       s>   	 �@     t       �>   	 #^A            �>    �jd     <1      �>   	 y0@     0       �>   	 jUA     �       �>   	 `�A     %       �>   	 @�A     �       �>     �f            �>   	 �N@     �       �>    �ae     �       �>   	 0j@            �>     [e            �>    �i            �>   	 �A     �      ?   	 �(B     *       ?    �Ze            '?   	 �@     �       :?   	 /CB            �A   	 ۲@     '       ]?   	 �R@     x       f?   	 t�A     %       v?   	 {$B     �       }?   	 n#B     �       �?    �6f            �                     �?   	 ��A            �?   	 :�A     
       �?   	 H�@     e      �?   	 �)B     �       �?   	 ��@     D       �?    `�g            �?   	 �@     m       �?   	 �]@     �      @   	 3�@            @   	 �1@            @   	 �A     �       /@   	 ��@            ;@   	 �.B            P@    �Pe            �/                     _@   	 Ӎ@            i@   	 �cA     !       r@    �f            z@   	 �/A     [       �@   	 �{A            �@   	 7�@     _       �@    (Re            �@   	 �A     �       �@   	 UvA            �@   	 Һ@            �&    @]d     0       �@   	 ��@     	      �@    ԓe            �@   	 ��@     R       A   	 �|A     -       A   	 �A     �       0A   	 �B     �       :A     Ze     �       CA   	 ��A     %       LA   	 &�A            XA    �6f            dA   	 �E@     �       uA    �if            �A    �Te     �       �A   	 �@     �       �A   	 Q�@     '       �A    Wf            �A    �i            �A   	 �HB             �A   	 �5B     Q       �A   	 O@     F       �A   	 ��@     $      B    ؓe             B    $�f            B   	 �hA     k       0B     �f            <B   	 I�@     I       IB    @Qe            [B   	 ��A     �       lB   	 �B     �       wB    @�f      @      �B   	 �@     U       �B   	 [�@     M       �B   	 �A     �       �B    �Qe            �B   	 ��A     �      �B    Ef            �B    Re            �B    @g            �B    �7e            C   	 ��@     `      C   	 .QA     p       C    �Jf            #C    ��e     H       0C    `g     �      @C   	 ��A     �       TC   	 ��@     
       eC   	 %@     �       rC    �i            {C     .f            �C   	 �A            �C   	 "A     �       �C   	 �f@     A       �C   	 �0B     &       �C   	 +�A     #       �C   	 ΍@            �C    Re            �C    x9f            �C    P`f            D    ��B            D    H�i            D    `Re             D    ��e            �    X`f            )D   	 ��@     Q       7D   	 ��@     �      ID    H_f            UD   	 6�A     B      iD   	 �@     (       �    �9f            tD   	 ��@     �       �D    �9f            �D   	 OB     �      >    ``f            �D   	  �@            �D   	 ��A           �D   	 Ƕ@     >       �D                     �D    ,Re            �D    �9f            �D    h�f            �D   	 f�A           E    �if            E   	 ��@             E   	 �3A     ,       !E   	 8A     �       6E   	 �A            BE    Ef            JE   	 ��@     "       TE   	 ߇@            dE    Ef            rE     Ef            ~E   	 _O@     �       �E     �i     P       �E    �Jf            �E   	 xB     ?       �E    h`f            �E    �`f            �E    �g            �E   	 h�@     Q       �E   	 ��@            �E    �Xe     �       F    Qe            F   	 ?A     
       &F    p�e            2F    (�f            =F   	 ^@     ^       JF   	 ��@     I       WF    �dd     �       ]F   	 t�@     �       uF   	 ��@            �F   	 x�@     �      �F   	 }�A     �      �F    �Pe            G    ��g     �      �F    �Qe            �F   	 �*A     2       �F   	 G@     u       �F    `^e     4      �F    �;f            �F    ��e            G    L�i            G   	 v�@     "       G    p�i            #G   	 ҹA            1G   	 #�A     �       KG   	 7�@     
       WG    `jd             dG    �;f            jG    �4g            tG   	 ee@     �       �G    �4g            �G    P�i            �G   	 �T@     )       �G   	 �@     �      �G   	 -@             �G                     �G   	 .@     �       �G   	 �@            �G   	 `A     �       H   	 A�A            H   	 Q@     V       'H    �6f            2H   	 ��@     "       FH   	 �C@     t       XH   	 fu@     D      jH   	 �QA     C      uH    0�f            �H   	 qB     �       �H   	 �'@            �H   	 �cA     4       �H    �Se     (       �H   	 VA     �      �H   	 و@            �H   	 -'@     �       �H   	 ��A     n       I   	 ��@     �       I   	 ��@     =       %I    ��e            7I   	 ��A            DI    �6f            NI   	 �1A     ?       [I    �jf            cI  " 	 �DB     �       rI  " 	  JB            yI   	 ��@           �I    �Pe            �I   	 әA     �       �I   	 �(A     -       �I   	 �@     �       �I   	 �?B           �I   	 ��@     
       �I   	 &�A     �      J   	 �f@            J   	 R�A     &       "J   	 �
B     �       5J   	 �B     9      IJ     _d     @       VJ   	 KA     d      hJ   	 H�@     n       tJ    �jf      @      }J   	 E!B     )       �J    0_f            �J   	 �@     $       �J   	 n�A     /       �J   	 �D@            �J    @^f     �       �J   	 ��@            C>    @Ye     �       ("     5g      @      �J   	 �e@     �       �J   	 e�A            �J   	 a9@     �       �J   	 "�A     �       K   	 �{@     l        K    (Ef            1K    �Qe            JK   	 ��@     �       [K   	 �/@            sK   	 ��@     u       �K    �;f            �K   	 u�A     �       �K    Qe            �K   	 �@            �K    `Ve            �K   	 ��A            �K   	 ��@     �       �K    0Ef            �K   	 Nq@     �      L   	 S3A     .       L   	 Ƈ@            $L    ��f            )L    T�i            1L   	 ��A     �       >L   	 5�@     &       RL   	 �V@     �       bL   	 G~@            �=    8�f            rL    @�f            �L   	 �yA     �      �L    �^d            �L   	 �=B            �L   	 	+A     <       �L    H�f            �L   	 �A     5      �L    ��i            �L    Ȫf            
M   	 �QA     W       !M   	 �B            .M   	 �t@     �       ?M   	 ��A     �       KM     �e     H       WM   	 �A     �      gM    �Qe            sM   	 WF@           �M   	 �i@     4       �M   	 ��@            �M    �Pe            �M   	 ?�@     8      �M   	 &@     !       �M   	 �A     �       �M    @Hf            �M    �ed            �M   	 pcA     2       �M    p�f            �M    DHf            N   	 [�@     �       N   	 s�@     d       'N    �Jf            .N   	 ?jA     _      ?N  " 	 �IB            FN   	 ��A     T       _N   	 ��A             mN   	 �*@            {N   	 '�@            �N    �%f            �N    $.f            �N    l`f            �N    p`f            �N  " 	 �IB     )       �N    P�f            �N    @3e     X      �N    P_f            �N   	 �o@     ?       �N   	 \4A     �       �N  " 	 �EB     -       	O    �Qe            O   	 3A            $O    LRe            -O   	 ��A     {      >O  " 	  FB     �       ZO    �Jf            `O   	 ��A     K       kO   	 }�A            {O   	 �c@     �      �O    X�i            �O   	 }�@     n       �O    �Jf            �O    t�f            �O   	 ��A     B       �O    �cf            �O    x�f            �O   	 ��A            �O     Bf     �      �O   	 ��A     �        P   	 �@     6       P    |�f            P   	 x�A     Z      %P   	 ,�@     y       1P   	 ע@     =       ;P   	 8-B            NP    �cf            ^P    @�e     H       vP   	 �'B     q       �P   	 �?B     0       �P    ��e     H       �P   	 )B     
       �P   	 n!B     f       �P   	 �A     �      �P   	 o�A           �P   	 ��A     �       �P                     �P   	 q�@            �P   	 Q�@            Q    �;f            Q    �;f            Q   	 �A     s       1Q   	 �}@            HQ   	 Q�@     )       SQ   	 ]�@     V       `Q   	 f�@     �       lQ    �ed            �Q    �Jf            �Q    HEf            �Q    \�i            �Q   	 �T@            �Q   	 e�@     .       �Q    �Qe            �Q     �e     H       �Q     �g            �Q    �Jf            �Q    X�f            �Q     �g      L     R    Гe            R   	 i�@     7       R   	 �B     �       3R                     AR                     GR   	 ]�A     D       PR    �,f     |       [R   	 p�@     �      nR    �Jf            xR   	 �@     4       h                      �R    4_f            �R   	 Q�A     �       �R   	 ��@            �R   	 �.B            E    x`f            �R    (.f            �R   	 yB            �R   	 ��@     �       �R   	 �@           �R    ��f            S     �h            
S    @�h            S    8_f            S   	 ��@     
       ,S    DRe            <S    ��f            KS     [e             RS    X-f            [S                     cS    �;f            oS    �`f            zS   	 X-A     E       �S    `�i            �S     Wf            �S   	 ˥@     ,       �S   	 B     �      �S   	 �@            �S    ,.f            �S    �Jf            y    `Hf            �S    ��f            �S    Df            T   	 �b@     �       T   	 u�A           T   	 4�@     2       *T   ؓe             6T   	 �@     �       =T   	 ��A     )       GT    �Pe            YT    0.f            eT   	 �@     &       mT    PEf            {T    XEf            �T    \-f            �T    ��e            �T    d�i            �T    �Pe            �T   	 +�@     <       �T    �Te     (       �T   	 �.B            �T    8Qe            �T   	 �,@            �0    ��f            �T   	 �"B     �       U    h�i            U   	 ��@            %U    �;f            -U   	 +�A            :U    4.f            BU   	 ��@     7       MU    @.f            TU   	 h�@     #       cU                     hU   	 ��@            rU   	 ۀ@     �      |U   	 �J@     �      �U   	 �dA     8       �U   	 �B     _       �U   	 R-B            �U   	 )B     2       �U   	 A     G       �U   	 ��@     h       �U   	 %�@            �U    ��f            �U    ��f            V    @[e     $       V    8(f            V  " 	 vEB            #X    �^d     p       'V   	 �@     y      :V   	 LvA     	       JV    `Ef     �       ZV   	 x�A     }      jV    (�i            sV   	 �S@     4      V                     �V   	 }5A     &       �V   	 �@     �       �V   	 *�@     A       �V    lQe            �V   	 N�@     V       �V    �7e            �V                     �V   	 'A     �       �V    �;f            W  " 	 �EB     -       W   	 oJ@     �       'W   	 @     N       9W   	 eD@     3       LW    �Qe            ^W    �;f            hW   	 N�A     -       |W   	 \[A     �      �W   	 ��@     
       �W   	 f�@     �      �W    xif            �W   	 jA     �       �W    �`f            �W    Qe            �W                     �W   	 h�A     �       �W   	 ��@     E       �W   	 C�@     H      X   	 ��A     �       X    H�h            X    �]d            0X   	 A     �      @X    ��e            NX    `Ff     �       XX   	 �7@            eX   	 S-B            pX    �Jf            �X   	 ,>A     �       K     -f            �X    Re            �X   	 v�A     �       �X   	 :�A     :       �X   	 �A     �       �X    �;f            �X   	 �3A     �       �X   	 �V@     U       �X    ؓe             �X    l�i            Y   	 �A     ,       Y     ug           Y    �e            'Y   	 ��@     �      6Y   	 �A            EY   	 ��A            PY   	 ��@     %       aY   	 �@     �       lY   	 �DB     &       �Y   	 �7A     �       �c    x�i            �Y   	 	�@     "      �Y   	 ��@     :       �Y   	 �A     p      �Y    zg            �Y    p�i            �Y   	 j2B     �        Z   	 �B     r       Z   	 )�@     �      Z   	 ?B     D       @Z   	 ��A     �       GZ    zg            BR                     SZ    \Qe            bZ   	 ��A     �       qZ    �6f            Z   	 �xA     �       �Z   	 �BB     �       �Z   	 ��A     f       �Z    H-f            �Z                     �Z   	 F1B     D       �Z   	 ��@     �        [    0�i            [    P�h            [  " 	 ;JB            "[   	 �'A     �       /[    �gf     �      :[   	 z�@            F[     Gf            P[   	 �k@            a[   	 $�@            n[   	 S=A     �       �[     �e     H       �[   	 y�A     �       �[   	 +AB     �       �[    X�h            �[   	 v�A     �       �[   	 --@     �      �[    �Qe            �[    P�e            �[   	 :A     Y       \    �;f            \   	 �y@            &\    �`f            1\   	 ��@     n       E\   	 M�@           R\    zg            \\    `�f            m\    �`f            y\   	 a�@     @       �\    @2f            �\   	 �}@            �\    ��f            �\   	 �5B     J      �\   	 �@            �\   	 �	A     X       �\   	 �A     !      ]    t�i             ]    ��i            -]   	 g�@     `       6]   	 K�@     Q       @]     Yf            O]   	 ��@           V]   	 ,�@     R       d]   	 �HB             z]    zg            �]    0Re            �]    �Qe            �]   	 *,@     �       �]    h�f            �]   	 �m@     �       �]    h6f            �]    ȓe            �]    �Pe            �]    �Jf            �]    zg            �]    x�i            ^   	 w�@     u       ^    �Jf            (^   	 �A     �      9^    Ъf            A^    |�i            L^    zg            R^   	 �n@     �       _^    �Pe            r^   	 �y@            }^   	 [5@     �       �^   	 ��@            �^    D2f            �^   	 `:@     =	      �^    XRe            �^    �Pe            �^   	 ��A     j       �^    ��i     P       �^    �;f            �^    (Qe            �3    `2f            �^   	 J
B            _    0(f            _    p�f            X    8�i             _   	 *@     %       ,_   	 �@     W      9_   	 f@     E      J_     Kf     �      U_    �Jf            ]_    ��e            l_   	 �+B     �      {_    T_f            �_   	 �
B     6       �_                     �_    ��i            �_    Qe            �_   	 �XA     �       �_  " 	 �FB     "       �_   	 �!@     �       �_   	  �A           `  " 	 �FB     "       `   	 ��@            "    �[e            (`    �Vf            1`   	 ?A            C`   	 6�A     v       P`   	 �)@     k       _`    x�f            r`    �i            `   	 �@     �       �`   	 
:B     �      �`   	 ��@     f       �`    TQe            �`   	 R�@            �`     Af            �`   	 |�A            a   	 �@B     6       %a    ��f            5a   	 H�@     "       Ba   	 !B     &       Ra    Qe            `a   	 v�@     a       la   	 [�A     &       za   	 �/B     �       �a    ��i            �a   	 �B            �a   	 ��A     A       �a   	 �B     t       �a    �Ze            �a    `We     (       �a   	 ,7A     p       �a    �`f            �a   	 \B           b   	 ��@            b    Qe            "b    `�h            -b    Af            6b   	 p<B     ?      _b   	 �oA     ~       mb   	 joA     �       ~b    @�e     �      �b     zg            �b   	 Ս@     K       �b   	 |V@     %       �b   	 ?@     #       �b   	 � @             �b     ^f            �b   	 � B     �       �b    Af            c   	 =�@     �       c   	 ��A     �      $c    ��i            0c   	 �.B            �    �Vf            :c    ��f            Lc   	 "�@            ]c   	 &B     \      gc   	 �DA     �       vc    �[e     �      c   	 :A     [       �c   	 ��@     -       �c   	  �@     
       �c   	 �@           �c   	 �@     �      �c   	 ��@            �c   	 
B     #       �c    ��f            �c    `�e            �c   	 �B     �       d    ��i            d   	 ��@            'd                     -d   	 $�A     Z       9d    `6f            Ed   	 �B     k       Xd     Af     �       _d   	 2�@            jd    ��i            vd   	 7:@     )       �d                     �d    @Df             �d   	 6:@            �d   	 ��@     8       �d    ��h      �      �d   	 ԍ@            �d     �d     �      �d    ��f            0<    ��i     �      �d    ��f            �d   	 ��A     �       e    �Qe            e   	 T
A     �       'e   	 ל@     U       6e   	 �@     )       De     Ze             crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.5424 dtor_idx.5426 frame_dummy object.5436 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux i_main.c doomgeneric_lemon.cpp addKeyToQueue _ZL20s_KeyQueueWriteIndex _ZL10s_KeyQueue _ZL19s_KeyQueueReadIndex _GLOBAL__sub_I_window dummy.c am_map.c f_w scale_ftom f_h m_y2 m_x2 old_m_x old_m_y old_m_w old_m_h followplayer plr markpointnum markpoints min_y min_x max_y max_x max_h min_scale_mtof max_scale_mtof m_paninc f_oldloc amclock lightlev ftom_zoommul mtof_zoommul st_notify.5921 marknums f_y f_x st_notify.5954 lastlevel.5958 lastepisode.5959 bigstate.5970 buffer.5971 cheating nexttic.5982 litelevelscnt.5984 litelevels.5983 fuck.6022 fl.6029 l.6048 their_colors.6078 d_event.c eventhead events eventtail d_iwad.c DirIsFile BuildIWADDirList num_iwad_dirs iwads d_loop.c PlayersInGame local_playeringame GetAdjustedTime new_sync BuildNewTic maketic ticdata skiptics recvtic player_class oldentertics.3134 frameon oldnettics frameskip d_main.c D_Endoom oldgamestate.6256 borderdrawcount.6257 fullscreen.6255 inhelpscreensstate.6254 viewactivestate.6252 menuactivestate.6253 packs.6339 gameversions d_mode.c valid_modes valid_versions CSWTCH.5 d_net.c RunTic exitmsg.4882 doom_loop_interface f_finale.c textscreens laststage.5474 f_wipe.c wipe_scr wipe_scr_end wipe_scr_start go wipes.2734 g_game.c gamekeydown mousearray joyarray joyxmove turnheld joyymove joystrafemove dclicks next_weapon weapon_order_table weapon_keys dclickstate dclicktime dclickstate2 dclicktime2 dclicks2 savegameslot carry.7153 savedescription CSWTCH.372 CSWTCH.370 resultbuf.7446 turbomessage.7213 hu_lib.c hu_stuff.c headsupactive message_on w_message message_nottobefuckedwith w_title w_chat w_inputbuffer always_off message_counter chat_dest chatchars altdown.5463 num_nobrainers.5467 lastmessage.5460 i_endoom.c i_joystick.c usejoystick joystick_physical_buttons joystick_index joystick_x_axis joystick_y_axis joystick_strafe_axis joystick_x_invert joystick_y_invert joystick_strafe_invert i_sound.c sound_module music_module i_system.c exit_funcs already_quitting firsttime.3501 mem_dump_dos622 dos_mem_dump mem_dump_win98 mem_dump_dosbox mem_dump_custom i_timer.c basetime m_argv.c m_bbox.c m_cheat.c m_config.c SearchCollection GetDefaultForName doom_defaults extra_defaults ParseIntParameter default_main_config default_extra_config scantokey extra_defaults_list doom_defaults_list m_controls.c m_fixed.c m_menu.c detailNames msgNames y.6469 x.6468 joywait.6441 mousewait.6442 lasty.6444 mousey.6443 lastx.6446 mousex.6445 m_misc.c m_random.c rndtable p_ceilng.c p_doors.c p_enemy.c easy.6345 p_floor.c p_inter.c p_lights.c p_map.c baseaddr.6206 p_maputl.c InterceptsMemoryOverrun intercepts_overrun InterceptsOverrun.part.0 p_mobj.c dummy_mobj.5937 p_plats.c p_pspr.c DecreaseAmmo p_saveg.c saveg_write8 saveg_write16 saveg_write32 saveg_write_thinker_t saveg_write_ceiling_t saveg_write_pad saveg_read8 saveg_read16 saveg_read32 saveg_read_pad saveg_read_thinker_t filename.5741 filename.5745 filename_size.5746 p_setup.c null_sector_is_initialized.6448 null_sector.6449 totallines p_sight.c p_spec.c first.6424 tmp_s3_floorheight.6425 tmp_s3_floorpic.6426 p_switch.c p_telept.c p_tick.c p_user.c r_bsp.c r_data.c r_draw.c background_buffer r_main.c r_plane.c r_segs.c r_sky.c r_things.c cliptop clipbot sha1.c Transform statdump.c num_captured_stats st_lib.c st_stuff.c ST_loadCallback ST_loadUnloadGraphics tallnum shortnum tallpercent faceback sbar ST_unloadCallback st_statusbaron st_firsttime plyr buf.6266 oldhealth.6275 lastcalc.6274 priority.6283 st_faceindex st_facecount oldweaponsowned st_oldhealth lastattackdown.6282 st_randomnumber largeammo.6291 w_ready st_fragscount st_notdeathmatch st_armson st_fragson st_msgcounter st_clock st_palette lu_palette w_ammo w_maxammo w_health w_arms w_armor w_armsbg w_faces w_keyboxes w_frags st_oldchat st_stopped s_sound.c S_StopChannel S_AdjustSoundParams snd_SfxVolume mus_playing mus_paused tables.c v_video.c dest_screen patchclip_callback wi_stuff.c WI_loadCallback WI_loadUnloadData NUMCMAPS lnames wiminus wbs yah splat NUMANIMS anims epsd1animinfo finished entering sp_secret colon timepatch sucks killers victims total bp background WI_unloadCallback lnodes bcnt acceleratestage snl_pointeron plrs dm_state cnt_pause dm_frags dm_totals bstar ng_state cnt_frags cnt_secret cnt_items cnt_kills dofrags sp_state cnt_par cnt_time epsd0animinfo epsd2animinfo w_checksum.c num_open_wadfiles w_file.c w_main.c w_wad.c lumphash unique_lumps z_zone.c w_file_stdc.c W_StdC_CloseFile W_StdC_OpenFile i_input.c shiftdown shiftxform i_video.c colors s_Fb doomgeneric.c ipc.cpp graphics.cpp window.cpp ../src/gfx/sse2.asm memcpy_sse2.loop memcpy_sse2_unaligned.loop memset32_sse2.loop memset32_sse2.ret memset64_sse2.loop memset64_sse2.ret runtime.cpp dstrings.c info.c sounds.c i_cdmus.c i_scale.c memio.c doomstat.c d_items.c _DYNAMIC _GLOBAL_OFFSET_TABLE_ EV_DoFloor _ZN4ListIP6WidgetED2Ev gametic consoleplayer usegamma main WI_updateNoState messageRoutine P_InitPicAnims I_StartSound R_CheckBBox _Z18memset32_optimizedPvjm cacheddistance buttonlist EpiDef M_DrawSaveLoadBorder I_UpdateSoundParams key_fire joybstrafe M_ChangeMessages validcount SHA1_Update EV_DoPlat AM_Drawer joybspeed S_Init stderr P_FindMinSurroundingLight devparm spryscale P_RemoveActiveCeiling P_GiveCard secondslideline R_ScaleFromGlobalAngle bodyque net_client_connected messx I_PrintStartupBanner _Z19HandleMouseMovementP6Window8Vector2i WritePCXfile Z_DumpHeap M_TempFile STlib_initMultIcon PIT_StompThing lumpinfo joybmenu R_DrawSpan epi remove M_ClearMenus casttics P_TempSaveGameFile A_SPosAttack messy pspriteiscale P_CalcSwing G_PlayerFinishLevel R_CheckPlane AM_findMinMaxBoundaries HU_Start M_VerifyNightmare _ZN4ListIP6WidgetE9remove_atEj A_Fall clipammo V_DrawShadowedPatch finesine HU_Stop A_Light0 PIT_AddLineIntercepts S_SetMusicVolume P_SlideMove ReadMenu1 realloc S_StopSound STlib_initBinIcon A_Light2 viewsin transcolfunc key_weapon5 M_Random ds_colormap A_Light1 PIT_RadiusAttack numspritelumps WI_drawStats D_Display message_dontfuckwithme key_weapon3 memset64_sse2 key_weapon2 messageNeedsInput key_weapon1 netgame weaponinfo A_LoadShotgun2 A_Hoof timingdemo AM_addMark R_RenderSegLoop messageToPrint WI_updateDeathmatchStats M_QuickSaveResponse lastanim wipe_exitColorXForm _ZN4ListIP6WidgetED1Ev bombspot key_invend W_CacheLumpName D_SuggestIWADName P_SpawnFireFlicker numbraintargets key_lookdown G_CheckDemoStatus I_SetWindowTitle M_WriteFile P_FindSectorFromLineTag P_SetThingPosition tmymove inhelpscreens P_CheckAmmo cht_CheckCheat numsprites P_ActivateInStasisCeiling W_LumpNameHash P_UnArchiveThinkers G_CmdChecksum sscanf M_SaveSelect gamemission M_StopMessage P_LoadSideDefs key_menu_right R_AddPointToBox S_music P_LineAttack HUlib_eraseIText P_NightmareRespawn savename wipe_initMelt DG_SleepMs episodes_e P_HitSlideLine spanstop offsetms EV_LightTurnOn key_menu_endgame PTR_UseTraverse M_GetIntVariable key_menu_forward rw_normalangle A_TroopAttack A_Explode timelimit R_PointInSubsector NewGameMenu A_VileTarget AM_drawGrid testcontrols_mousespeed dc_colormap forwardmove SHA1_Final D_ValidGameMode WI_Start D_GrabMouseCallback messageLastMenuActive quitsounds key_invpop G_DoSaveGame M_StartMessage nomonsters secretexit A_SargAttack R_InitFlats finaleflat V_DrawBlock _fini M_StringConcat P_SetupPsprites AM_rotate finetangent _Z13_CreateWindowP10win_info_t _Z5floord myargc _ZN6WindowC1Ev wipe_shittyColMajorXform opentop worldbottom A_BrainSpit A_FireCGun tempstring Z_ClearZone numlinespecials _ZN10win_info_tC2Ev G_InitNew P_MovePlayer MainDef texturecompositesize A_Fire totalsecret joybstraferight I_InitInput _ZN6WindowD2Ev key_left G_DeferedPlayDemo cachedxstep _ZdlPvm key_weapon4 key_weapon7 ST_updateFaceWidget finaletext V_DrawPatchDirect strcmp key_weapon6 I_SetGrabMouseCallback M_DrawEmptyCell V_SetPatchClipCallback G_Responder vissprites P_AddActivePlat key_menu_left key_weapon8 ST_calcPainOffset P_ExplodeMissile dc_source SaveMenu A_PosAttack M_LoadSelect sightzstart G_InitPlayer screenheightarray strace HU_Responder texturecomposite numvertexes I_ReadScreen D_PopEvent _Z24CreateFramebufferSurface6FBInfoPv M_vsnprintf D_PageDrawer P_TraverseIntercepts P_LoadNodes skytexturemid EV_DoLockedDoor HUlib_resetIText S_ChangeMusic gameepisode R_DrawColumnInCache R_PointToAngle key_message_refresh M_NewGame EV_DoDonut LoadMenu A_Lower numswitches aimslope configdir respawnmonsters Z_FreeTags WI_Ticker deathmatchstarts P_CheckSight _Znwm R_SetViewSize vanilla_savegame_limit W_NumLumps memset32_sse2 P_AddThinker P_InterceptVector2 texturememory P_Ticker planezlight sscount corpsehit M_ChooseSkill joybfire G_WorldDone M_DrawEpisode S_Start _Z12DrawGradientiiii10RGBAColourS_P7Surface A_FireMissile AM_drawPlayers P_TouchSpecialThing numpatches FixedMul F_Responder M_ApplyPlatformDefaults negonearray F_BunnyScroll ST_loadGraphics tmy R_Subsector spritememory worldlow HUlib_initIText R_DrawColumnLow mousebfire R_GenerateComposite malloc cachedheight M_SetConfigFilenames crushchange DG_Init dc_yl loopcount topslope ptflags G_BeginRecording A_KeenDie cheat_amap snd_channels NetUpdate A_FirePlasma numsubsectors tmx yspeed WI_slamBackground dc_yh centerxfrac HUlib_initTextLine EV_DoDoor chat_on fuzzpos setsizeneeded W_OpenFile D_PostEvent P_CrossBSPNode P_DropWeapon Z_Malloc wipegamestate _Z14ReceiveMessageP13ipc_message_t fflush S_SetSfxVolume key_arti_teleportother saveSlot strncmp A_BFGsound HUlib_addCharToTextLine ceilingplane system chat_macros FixedDiv framecount myargv fuzzoffset F_CastDrawer key_up sendsave _Z13DestroyWindowP6Window R_FillBackScreen doom1_endmsg HUlib_eraseTextLine M_ReadSaveStrings key_menu_gamma I_VideoBuffer_FB _Z8DrawRect4Rect10RGBAColourP7Surface A_BrainAwake strcpy pixhighstep levelTimeCount I_GetSfxLumpNum thintriangle_guy P_BlockLinesIterator P_CheckMissileSpawn A_BFGSpray walllights P_UseSpecialLine mouse_threshold rw_centerangle key_strafeleft singletics EV_BuildStairs D_StartNetGame mousebstraferight strrchr centeryfrac A_FirePistol key_menu_activate spritename netdemo distscale P_ChangeSwitchTexture M_ReadThis2 PIT_VileCheck show_endoom F_StartFinale R_InitTextures HUlib_delCharFromTextLine braintargeton finecosine I_UpdateSound cheat_clev rw_stopx A_SpawnFly A_FatAttack2 D_DoAdvanceDemo tantoangle HUlib_addPrefixToIText _ZN4ListIP6WidgetE10get_lengthEv _Z11PointInRect4Rect8Vector2i I_StopSong M_FileLength A_FatAttack1 longtics P_CrossSpecialLine A_OpenShotgun2 load_e P_DamageMobj P_FindHighestCeilingSurrounding P_ArchivePlayers A_PainAttack vileobj A_BspiAttack bfgedition P_GiveAmmo DG_GetKey R_InitColormaps V_RestoreBuffer fclose A_ReFire specials_e DG_SetWindowTitle W_ReleaseLumpNum R_PointToDist M_FileExists P_SpawnDoorCloseIn30 STlib_updateMultIcon bottomfrac key_arti_poisonbag T_PlatRaise M_snprintf showMessages M_ClearBox D_BindVariables I_UpdateNoBlit F_TextWrite oldgamestate _Z20DrawGradientVertical4Rect10RGBAColourS0_P7Surface key_jump M_QuitResponse AM_drawThings gameaction key_nextweapon precache P_BlockThingsIterator getNextSector AM_activateNewScale strdup HU_dequeueChatChar P_PathTraverse P_NewChaseDir vanilla_demo_limit detailshift WI_drawOnLnode M_DrawReadThis1 demo_p I_InitTimidityConfig extralight P_CrossSubsector spritetopoffset P_RespawnSpecials main_e lastopening P_ZMovement __mlibc_entry D_GameMissionString I_GraphicsCheckCommandLine M_ChangeSensitivity R_InitSpriteLumps __DTOR_END__ key_speed M_StringDuplicate tmthing WI_unloadData AM_Start I_GetTime ReadDef1 ST_Init P_TryMove A_WeaponReady key_strafe itemOn I_StopSound Z_FreeMemory I_InitMusic ReadDef2 P_InitThinkers slidemo sfxVolume AM_drawCrosshair M_SetConfigDir A_Look screensaver_mode cheat_choppers WI_drawEL P_GunShot blockmaplump topfrac WI_drawPercent R_AddLine M_DoSave soundtarget Z_FileDumpHeap strstr key_invright earlyout P_DivlineSide WI_drawNoState AM_drawLineCharacter R_RenderMaskedSegRange _Z8DrawRectiiiihhhP7Surface snd_sfxdevice HU_queueChatChar key_menu_down gameversion G_BuildTiccmd M_Options attackrange singledemo vfprintf _ZN8ListNodeIP6WidgetEC1Ev dclick_use rw_angle1 G_Ticker key_map_south _ZN10win_info_tC1Ev key_map_west P_SaveGameFile S_StartSound setdetail whichSkull P_FindHighestFloorSurrounding V_DrawVertLine iquetail WI_drawTime AM_loadPics AM_saveScaleAndLoc t2y rename scaledviewwidth leveltime P_SetPsprite P_ChangeSector P_UnArchivePlayers V_LoadXlaTable openbottom HUlib_addLineToSText Z_Init M_FindResponseFile I_GetPaletteIndex tmceilingz G_DoNewGame S_MusicPlaying key_map_follow demobuffer R_PointToAngle2 M_QuitDOOM spanfunc t2x SHA1_UpdateInt32 read_e A_BrainScream texturecolumnofs joybjump playerstarts demosequence PIT_AddThingIntercepts _Z14_DestroyWindowPv deathmatch_p angleturn shootthing castnum EV_DoCeiling numspechit key_invdrop M_StringEndsWith G_SaveGame key_invuse TRACEANGLE T_StrobeFlash pagename A_StartFire WI_End D_GetNumEpisodes AM_restoreScaleAndLoc P_GroupLines snd_musicdevice activeceilings cmap_to_fb P_SetMobjState V_DrawRawScreen A_PainShootSkull key_invleft P_ArchiveThinkers HUlib_eraseSText viewcos cmap_to_rgb565 R_DrawViewBorder I_PauseSong iwadfile M_BindStrifeControls EV_Teleport maskedtexturecol R_InitPointToAngle snd_musiccmd numlumps key_map_east ReadMenu2 R_ClipSolidWallSegment totalkills R_ClipPassWallSegment key_map_maxzoom A_VileChase strchr STlib_drawNum strncasecmp V_Init I_BeginRead numlines P_FindNextHighestFloor F_CastPrint WI_drawAnimatedBack M_BindMapControls S_sfx startmap P_BulletSlope P_PointOnLineSide I_SetPalette tmbbox R_NewVisSprite I_InitJoystick wipe_doColorXForm P_SpawnSpecials D_FindIWAD I_Endoom D_SuggestGameName A_BossDeath totalitems autostart P_PlayerInSpecialSector I_FinishUpdate key_arti_all key_usehealth st_backing_screen key_arti_egg projection mousebnextweapon viewwindowy bestslideline mousebstrafeleft A_FatRaise D_AdvanceDemo A_BrainDie snd_samplerate M_GetFloatVariable I_ResumeSong cheat_ammo V_DrawBox mousebprevweapon I_Quit V_DrawAltTLPatch M_GetSaveGameDir SaveDef SlopeDiv _Z10surfacecpyP7SurfaceS0_8Vector2i P_LoadSectors _Z11PaintWindowP6Window P_SpawnPlayerMissile A_SkullAttack spriteoffset P_SpawnPlayer thinkercap skytexture ftell key_map_grid key_multi_msg P_SpawnMapThing rw_scalestep finalecount bodyqueslot dc_texturemid mousey I_UpdateJoystick usething _ZN4ListIP6WidgetE8add_backES1_ D_IdentifyVersion R_DrawMasked A_SkelFist G_ExitLevel demoend menuactive ST_refreshBackground _Z18memset64_optimizedPvmm P_AddActiveCeiling V_DrawTLPatch AM_maxOutWindowScale I_DisplayFPSDots numnodes Z_ChangeTag2 WI_fragSum key_menu_detail sidedef W_Read castorder R_RenderPlayerView M_BindVariable AM_changeWindowScale modifiedgame spanstart planeheight fwrite R_ExecuteSetViewSize ST_initData P_UnsetThingPosition DG_ScreenBuffer OptionsDef EV_CeilingCrushStop key_map_zoomout P_MakeDivline HUlib_keyInIText P_AproxDistance P_LookForPlayers I_EndRead ds_xfrac starttime mousebbackward R_InitData G_DoCompleted tmfloorz maxframe key_arti_blastradius pixlow ds_source P_SpawnMissile worldhigh key_use viewheight M_ReadFile WI_checkForAccelerate flatmemory ST_unloadData worldtop getSide key_menu_confirm I_GetTicks P_RemoveMobj M_LoadDefaults ST_doRefresh ylookup clipangle viewwindowx M_BindWeaponControls P_RunThinkers mceilingclip WI_initVariables displayplayer HU_Init strncpy A_HeadAttack newend P_Thrust intercept_p tmdropoffz I_BindSoundVariables screenSize castdeath key_lookup key_map_mark P_UnArchiveSpecials W_ReleaseLumpName bmaporgy P_CalcHeight HUlib_drawTextLine W_CacheLumpNum M_EndGameResponse bmaporgx M_StringHeight dscount mapnames newvissprite putchar HUlib_drawSText mousebjump HUlib_addMessageToSText G_TimeDemo numtextures S_PauseSound mousebuse sprtemp P_LoadSubsectors P_SpawnMobj xlatab R_DrawFuzzColumnLow mousebstrafe M_DrawMainMenu P_UnArchiveWorld options_e P_GivePower M_StrCaseStr P_Init mobjinfo D_ProcessEvents P_LoadThings R_VideoErase V_CopyRect numflats F_Ticker checkcoord G_LoadGame diags vissprite_p R_DrawPSprite Z_ChangeUser screenblocks AM_changeWindowLoc _Z13HandleMouseUpP6Window8Vector2i F_Drawer V_DrawHorizLine Z_Free W_CheckCorrectIWAD finalestage StatDump ST_unloadGraphics PTR_AimTraverse I_GetEvent M_DrawNewGame cachedystep M_StrToInt G_DoLoadLevel P_NoiseAlert D_PageTicker R_RenderBSPNode A_BabyMetal I_BindVideoVariables joybnextweapon I_WaitVBL twoSided centery P_BringUpWeapon R_ClearDrawSegs A_BruisAttack key_flycenter ST_doPaletteStuff P_AllocateThinker M_ClearRandom T_MovePlane fb_scaling A_SkelMissile R_ClearClipSegs R_DrawMaskedColumn WI_drawLF gammamsg ST_Start ST_loadData castonmelee D_ConnectNetGame frontsector SoundMenu M_DrawThermo M_DrawReadThis2 test sprtopscreen memcpy_sse2 _Z8DrawRectiiii10RGBAColourP7Surface AM_Ticker M_StringJoin __bss_start lastspritelump P_ShootSpecialLine fuzzcolfunc A_CPosRefire key_map_clearmark ST_updateWidgets WI_drawNum viewangletox P_SpawnGlowingLight T_Glow P_AimLineAttack key_mission V_DrawMouseSpeedBox saveCharIndex key_arti_health centerx snd_cachesize A_Tracer P_LoadVertexes tmflags cheat_noclip scalelightfixed R_DrawPlayerSprites M_FinishReadThis AM_drawMarks dirtybox storedemo STlib_updateNum P_MobjThinker G_SecretExitLevel DG_GetTicksMs STlib_initPercent I_Sleep key_lookcenter lowres_turn blockmap gammatable rw_x quitsounds2 detailLevel M_StringWidth PTR_ShootTraverse save_stream R_InstallSpriteLump M_LoadGame PTR_SlideTraverse d_episode WI_updateStats M_CheckParm R_DrawSpanLow M_StringCopy fread key_flydown consistancy viewimage R_InitTextureMapping solidsegs HU_Erase A_GunFlash P_PointOnDivlineSide V_UseBuffer sound_e P_TryWalk I_ShutdownMusic quickSaveSlot currentMenu F_CastResponder vsprsortedhead bestslidefrac WI_Drawer numsides bottomslope scalelight M_BindChatControls M_ForceUppercase EpisodeMenu key_menu_save P_WriteSaveGameEOF musicVolume firstpatch AM_getIslope A_SpidRefire cpars I_BindJoystickVariables I_SetMusicVolume P_KillMobj R_MapPlane key_menu_quit key_demo_quit P_ActivateInStasis AM_LevelInit alphSwitchList turbodetected testcontrols pixlowstep M_AddToBox mfloorclip R_InitSprites R_DrawTranslatedColumnLow A_VileStart player_names d_map linecount G_DeathMatchSpawnPlayer viewplayer bottomstep wipe_exitMelt I_GetMemoryValue D_InitNetGame calloc AM_doFollowPlayer I_RegisterSong P_RadiusAttack SHA1_UpdateString F_DrawPatchCol castframes M_QuickLoadResponse D_ValidEpisodeMap G_WriteDemoTiccmd P_LoadSegs textureheight WI_updateAnimatedBack D_TryFindWADByName P_FindLowestFloorSurrounding LoadDef P_LoadLineDefs I_PrintDivider D_FindWADByName R_GetColumn A_FatAttack3 T_LightFlash main_loop_started S_StartMusic caststate P_FireWeapon linedef _ZN6WindowC2Ev _ZdaPv P_CheckMissileRange joybstrafeleft R_PointOnSegSide P_SubstNullMobj M_DrawOptions _Z12CreateWindowP10win_info_t M_ReadThis ST_Responder G_ScreenShot R_TextureNumForName WI_drawShowNextLoc WI_drawNetgameStats doom2_endmsg P_ArchiveSpecials M_WriteText drawsegs W_LumpLength bulletslope A_CloseShotgun2 ST_Stop D_IsEpisodeMap activeplats A_Pain G_DoReborn R_InitTables D_SetGameDescription V_DrawPatchFlipped HUlib_initSText skullAnimCounter key_arti_invulnerability P_RecursiveSound D_RegisterLoopCallbacks M_ExtractFileBase mousex R_InitLightTables key_menu_load M_SaveDefaultsAlternate OptionsMenu ST_diffDraw M_BindHexenControls saveOldString G_DoPlayDemo A_Raise I_PrecacheSounds ds_p topstep R_DrawColumn M_GetExecutableName wipe_ScreenWipe HUlib_drawIText texturecolumnlump P_PlayerThink gamemode _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i EV_StopPlat textures_hashtable P_XYMovement sttminus backsector GetSectorAtNullAddress WI_Responder G_ReadDemoTiccmd R_MakeSpans cheat_mypos R_ProjectSprite key_invhome D_CheckNetGame G_DoWorldDone A_Metal key_menu_incscreen I_Error AM_clearMarks R_InitTranslationTables viletryx sidemove getSector dc_iscale viletryy A_VileAttack P_SpawnLightFlash shootz P_UpdateSpecials _ZdlPv R_CheckTextureNumForName STlib_initNum D_QuitNetGame cht_GetParam tinttable fastparm bmapwidth numsectors _Znam lastflat sprnames savegame_error G_VanillaVersionCode A_Saw _ZN4ListIP6WidgetEC2Ev key_invquery A_CheckReload key_down R_StoreWallRange _ZN4ListIP6WidgetE6get_atEj nofit V_MarkRect V_LoadTintTable G_CheckSpot maskedtexture P_SpawnDoorRaiseIn5Mins openrange ds_x2 R_FlatNumForName levelTimer ds_y STlib_init hu_font V_DrawXlaPatch AM_unloadPics ds_x1 R_InitSpriteDefs I_InitSound M_EndGame I_ShutdownGraphics linespeciallist cheat_commercial_noclip Z_CheckHeap _Z12_PaintWindowPvi cheat_god Z_ZoneSize W_ReadLump PIT_CheckLine R_DrawPlanes ST_drawWidgets mkdir I_ShutdownJoystick A_SpawnSound demorecording viewactive P_InterceptVector HUlib_delCharFromIText P_GiveBody A_FaceTarget M_QuickSave mapnames_commercial floatok saveStringEnter bottomtexture wipe_initColorXForm I_AtExit key_pause cheat_mus basexscale bombsource spritewidth visplanes mouse_acceleration M_SfxVol WI_initNetgameStats __mlibc_errno fputs StatCopy windowInfo M_BindBaseControls la_damage M_DrawSelCell swingx R_PointOnSide A_FireCrackle I_EnableLoadingDisk startepisode W_CloseFile P_SpawnStrobeFlash AM_drawFline translations yslope baseyscale swingy M_MakeDirectory key_straferight dc_translation xspeed lasttime tolower defdemoname bmapheight P_RemoveActivePlat markfloor itemrespawntime M_StartControlPanel WI_drawDeathmatchStats AM_clearFB respawnparm linetarget dc_x chat_char G_PlayerReborn R_DrawSprite M_SaveGame __TMC_END__ M_Init ST_Ticker key_menu_messages advancedemo AM_Stop messageString read_e2 ticdup key_menu_screenshot rw_distance joybprevweapon A_PainDie SoundDef I_CheckIsScreensaver key_menu_up D_StartGameLoop W_GenerateHashTable toptexture P_Random d_skill R_InitSkyMap pagetic M_MusicVol mapdir A_PlayerScream atof I_Tactile HU_Ticker F_CastTicker P_FindLowestCeilingSurrounding WI_initStats I_StartFrame W_StdC_Read P_UseLines M_DrawLoad I_ConsoleStdout ds_xstep ds_ystep opposite usemouse _ZN6WindowD1Ev M_BindMenuControls P_RemoveThinker savegamestrings R_PrecacheLevel mainzone wipe_doMelt free A_FireBFG M_SetVariable M_StringStartsWith key_map_north P_CheckMeleeRange snd_maxslicetime_ms toupper P_SpawnPuff demoplayback _ZN4ListIP6WidgetEC1Ev F_StartCast AM_updateLightLev D_ValidGameVersion key_arti_teleport nodrawers STlib_updatePercent P_SetupLevel A_XScream A_Chase onground P_BoxOnLineSide numsegs key_menu_volume atoi R_DrawTranslatedColumn I_PrintBanner T_MoveCeiling R_FindPlane lastvisplane cheat_player_arrow P_CheckPosition stdc_wad_file endstring D_StartTitle I_StartTic secondslidefrac P_ReadSaveGameHeader key_useartifact R_DrawFuzzColumn V_DrawFilledBox R_ClearPlanes sendpause A_Punch wipe_EndScreen _edata rw_offset SHA1_Init xtoviewangle prndindex PIT_CheckThing R_ClearSprites S_Shutdown M_GetStrVariable M_DrawSave _Z9AddWidgetP6WidgetP6Window A_FireShotgun2 EV_VerticalDoor T_FireFlicker P_TeleportMove viewangleoffset rw_midtexturemid _Z16memcpy_optimizedPvS_m WI_loadData T_VerticalDoor _Z13_CreateWindowP10win_info_tPPvS2_ R_Init basecolfunc key_map_zoomin S_UpdateSounds castattacking P_DeathThink _Z15HandleMouseDownP6Window8Vector2i R_InitBuffer gamedescription fopen _Z11SendMessagem13ipc_message_t T_MoveFloor screenvisible ceilingfunc _ZdaPvm P_SpawnBlood switchlist P_GiveArmor newgame_e G_DeferedInitNew M_ParmExists P_WriteSaveGameHeader cheat_ammonokey STlib_updateBinIcon _Z17SwapWindowBuffersP6Window floorfunc R_SetupFrame TryRunTics key_spy drone P_LineOpening levelstarttic HUlib_clearTextLine blocklinks EV_TurnTagLightsOff P_GiveWeapon setblocks texturewidthmask sightcounts EV_StartLightStrobing startskill HUlib_eraseLineFromIText dccount _Z15DrawBitmapImageiiiiPhP7Surface M_SaveDefaults P_ThingHeightClip R_DrawVisSprite rw_toptexturemid spritelights A_Scream M_Episode itemrespawnque P_Move M_SizeDisplay memcpy_sse2_unaligned viewx key_flyup mousebforward D_ReceiveTic lastpatch G_DoLoadGame netcmds vanilla_keyboard_mapping key_menu_qload bombdamage viewz rw_bottomtexturemid I_ZoneBase ceilingline R_GenerateLookup curline midtexture viewy G_RecordDemo key_menu_decscreen HUlib_init D_DoomLoop A_CPosAttack startloadgame D_DoomMain key_right joybuse R_AddSprites overflowsprite players key_menu_back WI_initNoState I_VideoBuffer colormaps D_SaveGameIWADName AM_Responder AM_initVariables intercepts tmxmove key_prevweapon I_InitGraphics savegamelength WI_updateShowNextLoc memcpy rw_scale key_menu_abort P_LoadBlockMap _ZN8ListNodeIP6WidgetEC2Ev AM_drawWalls V_DrawPatch _ZN4ListIP6WidgetEixEj M_SetupNextMenu lowfloor P_ReadSaveGameEOF V_ScreenShot D_FindAllIWADs texturetranslation pspritescale M_BindHereticControls _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface M_DrawSound key_map_toggle I_MusicIsPlaying gameskill R_InitPlanes _Z12UpdateWindowP6Window flattranslation A_SkelWhoosh W_GetNumForName key_menu_help M_QuickLoad S_ResumeSound DG_DrawFrame skyflatnum WI_updateNetgameStats ST_Drawer WI_initDeathmatchStats mouseSensitivity NewDef A_FireShotgun rejectmatrix W_Checksum I_GetTimeMS key_menu_qsave floorplane usergame _Z10surfacecpyP7SurfaceS0_8Vector2i4Rect P_StartButton P_InitSwitchList cheat_powerup fixedcolormap M_CheckParmWithArgs wipe_StartScreen AM_minOutWindowScale AM_drawMline iquehead W_CheckNumForName gamemap A_BrainExplode ST_createWidgets segtextured dg_Create translationtables I_UnRegisterSong W_AddFile P_ArchiveWorld animdefs P_MovePsprites HU_Drawer M_Sound M_StringReplace AM_clipMline I_SoundIsPlaying WI_initShowNextLoc firstspritelump automapactive WI_initAnimatedBack pixhigh A_BrainPain fseek S_StopMusic savegamedir W_ParseCommandLine wminfo I_PlaySong markceiling PrintGameVersion strcasecmp key_multi_msgplayer PrintDehackedBanners I_ShutdownSound openings I_InitTimer states firstflat ds_yfrac R_SortVisSprites key_invkey PIT_ChangeSector M_ChangeDetail A_CyberAttack skullName  .symtab .strtab .shstrtab .interp .hash .dynsym .dynstr .rela.dyn .rela.plt .init .text .fini .rodata .eh_frame .init_array .ctors .dtors .dynamic .got .got.plt .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_str .debug_loc .debug_ranges .debug_macro                                                                               X@     X                                    #             h@     h      P                           )             �@     �      8                          1             �@     �      6                             9             (@     (      0                            C      B       X@     X      �                          M             0@     0                                    H             @@     @      �                            S             �@     �      �;                            Y             �JB     �J                                   _             �JB     �J     �                             g             ��C     ��     d}                             q             0Yd     0Y                                  }             8Yd     8Y                                   �             HYd     HY                                   �             XYd     XY     �                           �             �Zd     �Z                                  �             �Zd     �Z     `                            �             @\d     @\     �7                             �             ��e     ؓ     X%                             �      0               ؓ     +                             �                      �     �                             �                      ��                                   �                      ��     ?�                            �                      �W     ��                             �                      �Q     M1                            �                      �                                        0               �     �                                                �j     A�                                                 @4     �                             ,                     S     ��                                                   �F      �      !   �                	                      �!     Ne                                                   �j!     9                             